library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library Hast;
use Hast.SimpleMemory.all;

entity Hast_IP is 
    port(
        \DataIn\: In std_logic_vector(31 downto 0);
        \DataOut\: Out std_logic_vector(31 downto 0);
        \CellIndex\: Out integer;
        \ReadEnable\: Out boolean;
        \WriteEnable\: Out boolean;
        \ReadsDone\: In boolean;
        \WritesDone\: In boolean;
        \MemberId\: In integer;
        \Reset\: In std_logic;
        \Started\: In boolean;
        \Finished\: Out boolean;
        \Clock\: In std_logic
    );
    -- Hast_IP ID: ac8b1abb29548b4c174a7586ecf89e1be665a88547878a1f85ae430add66e46d
    -- (Date and time removed for approval testing.)
    -- Generated by Hastlayer - hastlayer.com
end Hast_IP;

architecture Imp of Hast_IP is 
    -- This IP was generated by Hastlayer from .NET code to mimic the original logic. Note the following:
    -- * For each member (methods, functions) in .NET a state machine was generated. Each state machine's name corresponds to 
    --   the original member's name.
    -- * Inputs and outputs are passed between state machines as shared objects.
    -- * There are operations that take multiple clock cycles like interacting with the memory and long-running arithmetic operations 
    --   (modulo, division, multiplication). These are awaited in subsequent states but be aware that some states can take more 
    --   than one clock cycle to produce their output.
    -- * The ExternalInvocationProxy process dispatches invocations that were started from the outside to the state machines.
    -- * The InternalInvocationProxy processes dispatch invocations between state machines.

    -- Enum declarations start
    type \Hast.Samples.SampleAssembly.SimdOperation\ is (
        \Hast.Samples.SampleAssembly.SimdOperation Hast.Samples.SampleAssembly.SimdOperation::Add\, 
        \Hast.Samples.SampleAssembly.SimdOperation Hast.Samples.SampleAssembly.SimdOperation::Subtract\, 
        \Hast.Samples.SampleAssembly.SimdOperation Hast.Samples.SampleAssembly.SimdOperation::Multiply\, 
        \Hast.Samples.SampleAssembly.SimdOperation Hast.Samples.SampleAssembly.SimdOperation::Divide\);
    -- Enum declarations end


    -- Custom inter-dependent type declarations start
    type \unsigned32_Array\ is array (integer range <>) of unsigned(31 downto 0);
    type \Hast.Samples.SampleAssembly.NumberContainer\ is record 
        \IsNull\: boolean;
        \WasIncreased\: boolean;
        \Number\: unsigned(31 downto 0);
    end record;
    type \Hast.Samples.SampleAssembly.NumberContainer_Array\ is array (integer range <>) of \Hast.Samples.SampleAssembly.NumberContainer\;
    type \boolean_Array\ is array (integer range <>) of boolean;
    type \signed32_Array\ is array (integer range <>) of signed(31 downto 0);
    type \Hast.Samples.SampleAssembly.MemoryContainer\ is record 
        \IsNull\: boolean;
    end record;
    -- Custom inter-dependent type declarations end


    -- System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::input declarations start
    -- Shared (global) variables:
    shared Variable \System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::input\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::input declarations end


    -- System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32).0 declarations start
    -- State machine states:
    type \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._States\ is (
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_0\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_1\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_2\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_3\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_4\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_5\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_6\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_7\);
    -- Signals:
    Signal \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._Finished\: boolean := false;
    Signal \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._Started\: boolean := false;
    Signal \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.indexObject.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32).0 declarations end


    -- System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32).1 declarations start
    -- State machine states:
    type \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._States\ is (
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_0\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_1\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_2\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_3\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_4\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_5\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_6\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_7\);
    -- Signals:
    Signal \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._Finished\: boolean := false;
    Signal \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._Started\: boolean := false;
    Signal \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.indexObject.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32).1 declarations end


    -- System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32).2 declarations start
    -- State machine states:
    type \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._States\ is (
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_0\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_1\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_2\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_3\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_4\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_5\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_6\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_7\);
    -- Signals:
    Signal \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._Finished\: boolean := false;
    Signal \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._Started\: boolean := false;
    Signal \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.indexObject.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32).2 declarations end


    -- System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32).3 declarations start
    -- State machine states:
    type \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._States\ is (
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_0\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_1\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_2\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_3\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_4\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_5\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_6\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_7\);
    -- Signals:
    Signal \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._Finished\: boolean := false;
    Signal \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._Started\: boolean := false;
    Signal \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.indexObject.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32).3 declarations end


    -- System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32).4 declarations start
    -- State machine states:
    type \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._States\ is (
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_0\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_1\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_2\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_3\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_4\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_5\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_6\, 
        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_7\);
    -- Signals:
    Signal \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._Finished\: boolean := false;
    Signal \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._Started\: boolean := false;
    Signal \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.indexObject.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32).4 declarations end


    -- System.Void Hast.Samples.SampleAssembly.ParallelAlgorithm::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations start
    -- State machine states:
    type \ParallelAlgorithm::Run(SimpleMemory).0._States\ is (
        \ParallelAlgorithm::Run(SimpleMemory).0._State_0\, 
        \ParallelAlgorithm::Run(SimpleMemory).0._State_1\, 
        \ParallelAlgorithm::Run(SimpleMemory).0._State_2\, 
        \ParallelAlgorithm::Run(SimpleMemory).0._State_3\, 
        \ParallelAlgorithm::Run(SimpleMemory).0._State_4\, 
        \ParallelAlgorithm::Run(SimpleMemory).0._State_5\, 
        \ParallelAlgorithm::Run(SimpleMemory).0._State_6\, 
        \ParallelAlgorithm::Run(SimpleMemory).0._State_7\, 
        \ParallelAlgorithm::Run(SimpleMemory).0._State_8\, 
        \ParallelAlgorithm::Run(SimpleMemory).0._State_9\);
    -- Signals:
    Signal \ParallelAlgorithm::Run(SimpleMemory).0._Finished\: boolean := false;
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.SimpleMemory.ReadEnable\: boolean := false;
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.SimpleMemory.WriteEnable\: boolean := false;
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).indexObject.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.0\: boolean := false;
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).indexObject.parameter.Out.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.1\: boolean := false;
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).indexObject.parameter.Out.2\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.2\: boolean := false;
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).indexObject.parameter.Out.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.3\: boolean := false;
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).indexObject.parameter.Out.4\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.4\: boolean := false;
    Signal \ParallelAlgorithm::Run(SimpleMemory).0._Started\: boolean := false;
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Finished.0\: boolean := false;
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Finished.1\: boolean := false;
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Finished.2\: boolean := false;
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Finished.3\: boolean := false;
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Finished.4\: boolean := false;
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).return.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).return.2\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).return.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).return.4\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.Void Hast.Samples.SampleAssembly.ParallelAlgorithm::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations end


    -- System.Void Hast.Samples.SampleAssembly.ObjectOrientedShowcase::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations start
    -- State machine states:
    type \ObjectOrientedShowcase::Run(SimpleMemory).0._States\ is (
        \ObjectOrientedShowcase::Run(SimpleMemory).0._State_0\, 
        \ObjectOrientedShowcase::Run(SimpleMemory).0._State_1\, 
        \ObjectOrientedShowcase::Run(SimpleMemory).0._State_2\, 
        \ObjectOrientedShowcase::Run(SimpleMemory).0._State_3\, 
        \ObjectOrientedShowcase::Run(SimpleMemory).0._State_4\, 
        \ObjectOrientedShowcase::Run(SimpleMemory).0._State_5\, 
        \ObjectOrientedShowcase::Run(SimpleMemory).0._State_6\, 
        \ObjectOrientedShowcase::Run(SimpleMemory).0._State_7\, 
        \ObjectOrientedShowcase::Run(SimpleMemory).0._State_8\, 
        \ObjectOrientedShowcase::Run(SimpleMemory).0._State_9\, 
        \ObjectOrientedShowcase::Run(SimpleMemory).0._State_10\, 
        \ObjectOrientedShowcase::Run(SimpleMemory).0._State_11\, 
        \ObjectOrientedShowcase::Run(SimpleMemory).0._State_12\, 
        \ObjectOrientedShowcase::Run(SimpleMemory).0._State_13\, 
        \ObjectOrientedShowcase::Run(SimpleMemory).0._State_14\, 
        \ObjectOrientedShowcase::Run(SimpleMemory).0._State_15\, 
        \ObjectOrientedShowcase::Run(SimpleMemory).0._State_16\, 
        \ObjectOrientedShowcase::Run(SimpleMemory).0._State_17\, 
        \ObjectOrientedShowcase::Run(SimpleMemory).0._State_18\, 
        \ObjectOrientedShowcase::Run(SimpleMemory).0._State_19\, 
        \ObjectOrientedShowcase::Run(SimpleMemory).0._State_20\, 
        \ObjectOrientedShowcase::Run(SimpleMemory).0._State_21\, 
        \ObjectOrientedShowcase::Run(SimpleMemory).0._State_22\);
    -- Signals:
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0._Finished\: boolean := false;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.SimpleMemory.ReadEnable\: boolean := false;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.SimpleMemory.WriteEnable\: boolean := false;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::.ctor(SimpleMemory).this.parameter.Out.0\: \Hast.Samples.SampleAssembly.MemoryContainer\;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::.ctor(SimpleMemory)._Started.0\: boolean := false;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::GetInput().this.parameter.Out.0\: \Hast.Samples.SampleAssembly.MemoryContainer\;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::GetInput()._Started.0\: boolean := false;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor().this.parameter.Out.0\: \Hast.Samples.SampleAssembly.NumberContainer\;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor()._Started.0\: boolean := false;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor(UInt32).this.parameter.Out.0\: \Hast.Samples.SampleAssembly.NumberContainer\;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor(UInt32).number.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor(UInt32)._Started.0\: boolean := false;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::set_NumberPlusFive(UInt32).this.parameter.Out.0\: \Hast.Samples.SampleAssembly.NumberContainer\;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::set_NumberPlusFive(UInt32).value.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::set_NumberPlusFive(UInt32)._Started.0\: boolean := false;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32).this.parameter.Out.0\: \Hast.Samples.SampleAssembly.NumberContainer\;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32).increaseBy.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32)._Started.0\: boolean := false;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::get_NumberPlusFive().this.parameter.Out.0\: \Hast.Samples.SampleAssembly.NumberContainer\;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::get_NumberPlusFive()._Started.0\: boolean := false;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).numberContainers.parameter.Out.0\: \Hast.Samples.SampleAssembly.NumberContainer_Array\(0 to 3);
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[])._Started.0\: boolean := false;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0._Started\: boolean := false;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::.ctor(SimpleMemory).this.parameter.In.0\: \Hast.Samples.SampleAssembly.MemoryContainer\;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::.ctor(SimpleMemory)._Finished.0\: boolean := false;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::GetInput().this.parameter.In.0\: \Hast.Samples.SampleAssembly.MemoryContainer\;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::GetInput()._Finished.0\: boolean := false;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::GetInput().return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor().this.parameter.In.0\: \Hast.Samples.SampleAssembly.NumberContainer\;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor()._Finished.0\: boolean := false;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor(UInt32).this.parameter.In.0\: \Hast.Samples.SampleAssembly.NumberContainer\;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor(UInt32)._Finished.0\: boolean := false;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::set_NumberPlusFive(UInt32).this.parameter.In.0\: \Hast.Samples.SampleAssembly.NumberContainer\;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::set_NumberPlusFive(UInt32)._Finished.0\: boolean := false;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32).this.parameter.In.0\: \Hast.Samples.SampleAssembly.NumberContainer\;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32)._Finished.0\: boolean := false;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::get_NumberPlusFive().this.parameter.In.0\: \Hast.Samples.SampleAssembly.NumberContainer\;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::get_NumberPlusFive()._Finished.0\: boolean := false;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::get_NumberPlusFive().return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).numberContainers.parameter.In.0\: \Hast.Samples.SampleAssembly.NumberContainer_Array\(0 to 3);
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[])._Finished.0\: boolean := false;
    Signal \ObjectOrientedShowcase::Run(SimpleMemory).0.ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.Void Hast.Samples.SampleAssembly.ObjectOrientedShowcase::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations end


    -- System.UInt32 Hast.Samples.SampleAssembly.ObjectOrientedShowcase::SumNumberCointainers(Hast.Samples.SampleAssembly.NumberContainer[]).0 declarations start
    -- State machine states:
    type \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._States\ is (
        \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State_0\, 
        \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State_1\, 
        \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State_2\, 
        \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State_3\, 
        \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State_4\);
    -- Signals:
    Signal \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._Finished\: boolean := false;
    Signal \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.numberContainers.parameter.Out\: \Hast.Samples.SampleAssembly.NumberContainer_Array\(0 to 3);
    Signal \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._Started\: boolean := false;
    Signal \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.numberContainers.parameter.In\: \Hast.Samples.SampleAssembly.NumberContainer_Array\(0 to 3);
    -- System.UInt32 Hast.Samples.SampleAssembly.ObjectOrientedShowcase::SumNumberCointainers(Hast.Samples.SampleAssembly.NumberContainer[]).0 declarations end


    -- System.Void Hast.Samples.SampleAssembly.NumberContainer::.ctor().0 declarations start
    -- State machine states:
    type \NumberContainer::.ctor().0._States\ is (
        \NumberContainer::.ctor().0._State_0\, 
        \NumberContainer::.ctor().0._State_1\, 
        \NumberContainer::.ctor().0._State_2\);
    -- Signals:
    Signal \NumberContainer::.ctor().0._Finished\: boolean := false;
    Signal \NumberContainer::.ctor().0.this.parameter.Out\: \Hast.Samples.SampleAssembly.NumberContainer\;
    Signal \NumberContainer::.ctor().0._Started\: boolean := false;
    Signal \NumberContainer::.ctor().0.this.parameter.In\: \Hast.Samples.SampleAssembly.NumberContainer\;
    -- System.Void Hast.Samples.SampleAssembly.NumberContainer::.ctor().0 declarations end


    -- System.Void Hast.Samples.SampleAssembly.NumberContainer::.ctor(System.UInt32).0 declarations start
    -- State machine states:
    type \NumberContainer::.ctor(UInt32).0._States\ is (
        \NumberContainer::.ctor(UInt32).0._State_0\, 
        \NumberContainer::.ctor(UInt32).0._State_1\, 
        \NumberContainer::.ctor(UInt32).0._State_2\);
    -- Signals:
    Signal \NumberContainer::.ctor(UInt32).0._Finished\: boolean := false;
    Signal \NumberContainer::.ctor(UInt32).0.this.parameter.Out\: \Hast.Samples.SampleAssembly.NumberContainer\;
    Signal \NumberContainer::.ctor(UInt32).0._Started\: boolean := false;
    Signal \NumberContainer::.ctor(UInt32).0.this.parameter.In\: \Hast.Samples.SampleAssembly.NumberContainer\;
    Signal \NumberContainer::.ctor(UInt32).0.number.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.Void Hast.Samples.SampleAssembly.NumberContainer::.ctor(System.UInt32).0 declarations end


    -- System.UInt32 Hast.Samples.SampleAssembly.NumberContainer::IncreaseNumber(System.UInt32).0 declarations start
    -- State machine states:
    type \NumberContainer::IncreaseNumber(UInt32).0._States\ is (
        \NumberContainer::IncreaseNumber(UInt32).0._State_0\, 
        \NumberContainer::IncreaseNumber(UInt32).0._State_1\, 
        \NumberContainer::IncreaseNumber(UInt32).0._State_2\);
    -- Signals:
    Signal \NumberContainer::IncreaseNumber(UInt32).0._Finished\: boolean := false;
    Signal \NumberContainer::IncreaseNumber(UInt32).0.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \NumberContainer::IncreaseNumber(UInt32).0.this.parameter.Out\: \Hast.Samples.SampleAssembly.NumberContainer\;
    Signal \NumberContainer::IncreaseNumber(UInt32).0._Started\: boolean := false;
    Signal \NumberContainer::IncreaseNumber(UInt32).0.this.parameter.In\: \Hast.Samples.SampleAssembly.NumberContainer\;
    Signal \NumberContainer::IncreaseNumber(UInt32).0.increaseBy.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.UInt32 Hast.Samples.SampleAssembly.NumberContainer::IncreaseNumber(System.UInt32).0 declarations end


    -- System.UInt32 Hast.Samples.SampleAssembly.NumberContainer::get_NumberPlusFive().0 declarations start
    -- State machine states:
    type \NumberContainer::get_NumberPlusFive().0._States\ is (
        \NumberContainer::get_NumberPlusFive().0._State_0\, 
        \NumberContainer::get_NumberPlusFive().0._State_1\, 
        \NumberContainer::get_NumberPlusFive().0._State_2\);
    -- Signals:
    Signal \NumberContainer::get_NumberPlusFive().0._Finished\: boolean := false;
    Signal \NumberContainer::get_NumberPlusFive().0.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \NumberContainer::get_NumberPlusFive().0.this.parameter.Out\: \Hast.Samples.SampleAssembly.NumberContainer\;
    Signal \NumberContainer::get_NumberPlusFive().0._Started\: boolean := false;
    Signal \NumberContainer::get_NumberPlusFive().0.this.parameter.In\: \Hast.Samples.SampleAssembly.NumberContainer\;
    -- System.UInt32 Hast.Samples.SampleAssembly.NumberContainer::get_NumberPlusFive().0 declarations end


    -- System.Void Hast.Samples.SampleAssembly.NumberContainer::set_NumberPlusFive(System.UInt32).0 declarations start
    -- State machine states:
    type \NumberContainer::set_NumberPlusFive(UInt32).0._States\ is (
        \NumberContainer::set_NumberPlusFive(UInt32).0._State_0\, 
        \NumberContainer::set_NumberPlusFive(UInt32).0._State_1\, 
        \NumberContainer::set_NumberPlusFive(UInt32).0._State_2\);
    -- Signals:
    Signal \NumberContainer::set_NumberPlusFive(UInt32).0._Finished\: boolean := false;
    Signal \NumberContainer::set_NumberPlusFive(UInt32).0.this.parameter.Out\: \Hast.Samples.SampleAssembly.NumberContainer\;
    Signal \NumberContainer::set_NumberPlusFive(UInt32).0._Started\: boolean := false;
    Signal \NumberContainer::set_NumberPlusFive(UInt32).0.this.parameter.In\: \Hast.Samples.SampleAssembly.NumberContainer\;
    Signal \NumberContainer::set_NumberPlusFive(UInt32).0.value.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.Void Hast.Samples.SampleAssembly.NumberContainer::set_NumberPlusFive(System.UInt32).0 declarations end


    -- System.Void Hast.Samples.SampleAssembly.MemoryContainer::.ctor(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations start
    -- State machine states:
    type \MemoryContainer::.ctor(SimpleMemory).0._States\ is (
        \MemoryContainer::.ctor(SimpleMemory).0._State_0\, 
        \MemoryContainer::.ctor(SimpleMemory).0._State_1\, 
        \MemoryContainer::.ctor(SimpleMemory).0._State_2\);
    -- Signals:
    Signal \MemoryContainer::.ctor(SimpleMemory).0._Finished\: boolean := false;
    Signal \MemoryContainer::.ctor(SimpleMemory).0.this.parameter.Out\: \Hast.Samples.SampleAssembly.MemoryContainer\;
    Signal \MemoryContainer::.ctor(SimpleMemory).0._Started\: boolean := false;
    Signal \MemoryContainer::.ctor(SimpleMemory).0.this.parameter.In\: \Hast.Samples.SampleAssembly.MemoryContainer\;
    -- System.Void Hast.Samples.SampleAssembly.MemoryContainer::.ctor(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations end


    -- System.UInt32 Hast.Samples.SampleAssembly.MemoryContainer::GetInput().0 declarations start
    -- State machine states:
    type \MemoryContainer::GetInput().0._States\ is (
        \MemoryContainer::GetInput().0._State_0\, 
        \MemoryContainer::GetInput().0._State_1\, 
        \MemoryContainer::GetInput().0._State_2\, 
        \MemoryContainer::GetInput().0._State_3\);
    -- Signals:
    Signal \MemoryContainer::GetInput().0._Finished\: boolean := false;
    Signal \MemoryContainer::GetInput().0.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \MemoryContainer::GetInput().0.this.parameter.Out\: \Hast.Samples.SampleAssembly.MemoryContainer\;
    Signal \MemoryContainer::GetInput().0.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \MemoryContainer::GetInput().0.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \MemoryContainer::GetInput().0.SimpleMemory.ReadEnable\: boolean := false;
    Signal \MemoryContainer::GetInput().0.SimpleMemory.WriteEnable\: boolean := false;
    Signal \MemoryContainer::GetInput().0._Started\: boolean := false;
    Signal \MemoryContainer::GetInput().0.this.parameter.In\: \Hast.Samples.SampleAssembly.MemoryContainer\;
    -- System.UInt32 Hast.Samples.SampleAssembly.MemoryContainer::GetInput().0 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32).0 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.return\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.numberObject.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32).0 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32).1 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.return\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.numberObject.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32).1 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32).2 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.return\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.numberObject.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32).2 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32).3 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.return\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.numberObject.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32).3 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32).4 declarations start
    -- State machine states:
    type \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._States\ is (
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_0\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_1\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_2\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_3\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_4\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_5\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_6\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_7\, 
        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_8\);
    -- Signals:
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._Finished\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.return\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._Started\: boolean := false;
    Signal \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.numberObject.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32).4 declarations end


    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumber(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations start
    -- State machine states:
    type \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._States\ is (
        \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_0\, 
        \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_1\, 
        \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_2\, 
        \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_3\, 
        \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_4\, 
        \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_5\);
    -- Signals:
    Signal \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Finished\: boolean := false;
    Signal \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.ReadEnable\: boolean := false;
    Signal \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.WriteEnable\: boolean := false;
    Signal \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).number.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\: boolean := false;
    Signal \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Started\: boolean := false;
    Signal \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\: boolean := false;
    Signal \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).return.0\: boolean := false;
    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumber(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations end


    -- System.Threading.Tasks.Task Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberAsync(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations start
    -- State machine states:
    type \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._States\ is (
        \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_0\, 
        \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_1\, 
        \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_2\, 
        \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_3\);
    -- Signals:
    Signal \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._Finished\: boolean := false;
    Signal \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\: boolean := false;
    Signal \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._Started\: boolean := false;
    Signal \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\: boolean := false;
    -- System.Threading.Tasks.Task Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberAsync(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations end


    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ArePrimeNumbers(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations start
    -- State machine states:
    type \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._States\ is (
        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_0\, 
        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_1\, 
        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_2\, 
        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_3\, 
        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_4\, 
        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_5\, 
        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_6\, 
        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_7\, 
        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_8\);
    -- Signals:
    Signal \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._Finished\: boolean := false;
    Signal \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\: boolean := false;
    Signal \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\: boolean := false;
    Signal \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).number.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\: boolean := false;
    Signal \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._Started\: boolean := false;
    Signal \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\: boolean := false;
    Signal \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).return.0\: boolean := false;
    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ArePrimeNumbers(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations end


    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations start
    -- State machine states:
    type \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._States\ is (
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_0\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_1\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_2\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_3\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_4\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_5\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_6\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_7\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_8\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_9\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_10\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_11\, 
        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_12\);
    -- Signals:
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._Finished\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).numberObject.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.0\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).numberObject.parameter.Out.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.1\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).numberObject.parameter.Out.2\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.2\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).numberObject.parameter.Out.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.3\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).numberObject.parameter.Out.4\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.4\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._Started\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Finished.0\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Finished.1\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Finished.2\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Finished.3\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Finished.4\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).return.0\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).return.1\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).return.2\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).return.3\: boolean := false;
    Signal \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).return.4\: boolean := false;
    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberInternal(System.UInt32).0 declarations start
    -- State machine states:
    type \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._States\ is (
        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_0\, 
        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_1\, 
        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_2\, 
        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_3\, 
        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_4\, 
        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_5\, 
        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_6\, 
        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_7\, 
        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_8\);
    -- Signals:
    Signal \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Finished\: boolean := false;
    Signal \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.return\: boolean := false;
    Signal \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Started\: boolean := false;
    Signal \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.number.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberInternal(System.UInt32).0 declarations end


    -- System.Void Hast.Samples.SampleAssembly.RecursiveAlgorithms::CalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations start
    -- State machine states:
    type \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._States\ is (
        \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State_0\, 
        \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State_1\, 
        \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State_2\, 
        \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State_3\, 
        \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State_4\, 
        \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State_5\, 
        \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State_6\);
    -- Signals:
    Signal \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._Finished\: boolean := false;
    Signal \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.ReadEnable\: boolean := false;
    Signal \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.WriteEnable\: boolean := false;
    Signal \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\: boolean := false;
    Signal \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._Started\: boolean := false;
    Signal \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\: boolean := false;
    Signal \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.Void Hast.Samples.SampleAssembly.RecursiveAlgorithms::CalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations end


    -- System.Void Hast.Samples.SampleAssembly.RecursiveAlgorithms::CalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations start
    -- State machine states:
    type \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._States\ is (
        \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State_0\, 
        \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State_1\, 
        \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State_2\, 
        \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State_3\, 
        \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State_4\, 
        \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State_5\, 
        \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State_6\);
    -- Signals:
    Signal \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._Finished\: boolean := false;
    Signal \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.ReadEnable\: boolean := false;
    Signal \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.WriteEnable\: boolean := false;
    Signal \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\: boolean := false;
    Signal \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._Started\: boolean := false;
    Signal \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\: boolean := false;
    Signal \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.Void Hast.Samples.SampleAssembly.RecursiveAlgorithms::CalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).0 declarations start
    -- State machine states:
    type \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._States\ is (
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_0\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_1\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_2\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_3\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_4\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_5\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_6\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_7\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_8\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_9\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_10\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_11\);
    -- Signals:
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Finished\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.SimpleMemory.ReadEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.SimpleMemory.WriteEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Started\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.number.parameter.In\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).0 declarations end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).1 declarations start
    -- State machine states:
    type \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._States\ is (
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_0\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_1\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_2\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_3\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_4\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_5\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_6\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_7\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_8\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_9\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_10\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_11\);
    -- Signals:
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Finished\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.SimpleMemory.ReadEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.SimpleMemory.WriteEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Started\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.number.parameter.In\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).1 declarations end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).2 declarations start
    -- State machine states:
    type \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._States\ is (
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_0\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_1\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_2\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_3\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_4\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_5\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_6\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_7\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_8\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_9\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_10\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_11\);
    -- Signals:
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Finished\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.SimpleMemory.ReadEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.SimpleMemory.WriteEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Started\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.number.parameter.In\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).2 declarations end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).3 declarations start
    -- State machine states:
    type \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._States\ is (
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_0\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_1\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_2\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_3\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_4\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_5\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_6\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_7\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_8\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_9\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_10\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_11\);
    -- Signals:
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Finished\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.SimpleMemory.ReadEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.SimpleMemory.WriteEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Started\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.number.parameter.In\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).3 declarations end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).4 declarations start
    -- State machine states:
    type \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._States\ is (
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_0\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_1\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_2\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_3\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_4\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_5\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_6\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_7\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_8\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_9\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_10\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_11\);
    -- Signals:
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Finished\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.SimpleMemory.ReadEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.SimpleMemory.WriteEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Started\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.number.parameter.In\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).4 declarations end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).5 declarations start
    -- State machine states:
    type \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._States\ is (
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_0\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_1\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_2\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_3\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_4\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_5\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_6\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_7\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_8\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_9\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_10\, 
        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_11\);
    -- Signals:
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Finished\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.SimpleMemory.ReadEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.SimpleMemory.WriteEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Started\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.number.parameter.In\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).5 declarations end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).0 declarations start
    -- State machine states:
    type \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._States\ is (
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_0\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_1\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_2\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_3\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_4\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_5\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_6\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_7\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_8\);
    -- Signals:
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Finished\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.SimpleMemory.ReadEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.SimpleMemory.WriteEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Started\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.number.parameter.In\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).0 declarations end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).1 declarations start
    -- State machine states:
    type \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._States\ is (
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_0\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_1\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_2\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_3\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_4\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_5\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_6\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_7\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_8\);
    -- Signals:
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Finished\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.SimpleMemory.ReadEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.SimpleMemory.WriteEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Started\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.number.parameter.In\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).1 declarations end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).2 declarations start
    -- State machine states:
    type \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._States\ is (
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_0\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_1\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_2\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_3\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_4\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_5\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_6\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_7\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_8\);
    -- Signals:
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Finished\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.SimpleMemory.ReadEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.SimpleMemory.WriteEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Started\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.number.parameter.In\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).2 declarations end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).3 declarations start
    -- State machine states:
    type \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._States\ is (
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_0\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_1\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_2\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_3\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_4\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_5\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_6\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_7\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_8\);
    -- Signals:
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Finished\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.SimpleMemory.ReadEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.SimpleMemory.WriteEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Started\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.number.parameter.In\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).3 declarations end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).4 declarations start
    -- State machine states:
    type \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._States\ is (
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_0\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_1\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_2\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_3\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_4\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_5\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_6\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_7\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_8\);
    -- Signals:
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Finished\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.SimpleMemory.ReadEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.SimpleMemory.WriteEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Started\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.number.parameter.In\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).4 declarations end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).5 declarations start
    -- State machine states:
    type \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._States\ is (
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_0\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_1\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_2\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_3\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_4\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_5\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_6\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_7\, 
        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_8\);
    -- Signals:
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Finished\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.SimpleMemory.ReadEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.SimpleMemory.WriteEnable\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Started\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.number.parameter.In\: signed(15 downto 0) := to_signed(0, 16);
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\: boolean := false;
    Signal \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).5 declarations end


    -- System.Void Hast.Samples.SampleAssembly.SimdCalculator::AddVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations start
    -- State machine states:
    type \SimdCalculator::AddVectors(SimpleMemory).0._States\ is (
        \SimdCalculator::AddVectors(SimpleMemory).0._State_0\, 
        \SimdCalculator::AddVectors(SimpleMemory).0._State_1\, 
        \SimdCalculator::AddVectors(SimpleMemory).0._State_2\, 
        \SimdCalculator::AddVectors(SimpleMemory).0._State_3\);
    -- Signals:
    Signal \SimdCalculator::AddVectors(SimpleMemory).0._Finished\: boolean := false;
    Signal \SimdCalculator::AddVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).operation.parameter.Out.0\: \Hast.Samples.SampleAssembly.SimdOperation\;
    Signal \SimdCalculator::AddVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\: boolean := false;
    Signal \SimdCalculator::AddVectors(SimpleMemory).0._Started\: boolean := false;
    Signal \SimdCalculator::AddVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\: boolean := false;
    -- System.Void Hast.Samples.SampleAssembly.SimdCalculator::AddVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations end


    -- System.Void Hast.Samples.SampleAssembly.SimdCalculator::SubtractVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations start
    -- State machine states:
    type \SimdCalculator::SubtractVectors(SimpleMemory).0._States\ is (
        \SimdCalculator::SubtractVectors(SimpleMemory).0._State_0\, 
        \SimdCalculator::SubtractVectors(SimpleMemory).0._State_1\, 
        \SimdCalculator::SubtractVectors(SimpleMemory).0._State_2\, 
        \SimdCalculator::SubtractVectors(SimpleMemory).0._State_3\);
    -- Signals:
    Signal \SimdCalculator::SubtractVectors(SimpleMemory).0._Finished\: boolean := false;
    Signal \SimdCalculator::SubtractVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).operation.parameter.Out.0\: \Hast.Samples.SampleAssembly.SimdOperation\;
    Signal \SimdCalculator::SubtractVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\: boolean := false;
    Signal \SimdCalculator::SubtractVectors(SimpleMemory).0._Started\: boolean := false;
    Signal \SimdCalculator::SubtractVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\: boolean := false;
    -- System.Void Hast.Samples.SampleAssembly.SimdCalculator::SubtractVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations end


    -- System.Void Hast.Samples.SampleAssembly.SimdCalculator::MultiplyVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations start
    -- State machine states:
    type \SimdCalculator::MultiplyVectors(SimpleMemory).0._States\ is (
        \SimdCalculator::MultiplyVectors(SimpleMemory).0._State_0\, 
        \SimdCalculator::MultiplyVectors(SimpleMemory).0._State_1\, 
        \SimdCalculator::MultiplyVectors(SimpleMemory).0._State_2\, 
        \SimdCalculator::MultiplyVectors(SimpleMemory).0._State_3\);
    -- Signals:
    Signal \SimdCalculator::MultiplyVectors(SimpleMemory).0._Finished\: boolean := false;
    Signal \SimdCalculator::MultiplyVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).operation.parameter.Out.0\: \Hast.Samples.SampleAssembly.SimdOperation\;
    Signal \SimdCalculator::MultiplyVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\: boolean := false;
    Signal \SimdCalculator::MultiplyVectors(SimpleMemory).0._Started\: boolean := false;
    Signal \SimdCalculator::MultiplyVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\: boolean := false;
    -- System.Void Hast.Samples.SampleAssembly.SimdCalculator::MultiplyVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations end


    -- System.Void Hast.Samples.SampleAssembly.SimdCalculator::DivideVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations start
    -- State machine states:
    type \SimdCalculator::DivideVectors(SimpleMemory).0._States\ is (
        \SimdCalculator::DivideVectors(SimpleMemory).0._State_0\, 
        \SimdCalculator::DivideVectors(SimpleMemory).0._State_1\, 
        \SimdCalculator::DivideVectors(SimpleMemory).0._State_2\, 
        \SimdCalculator::DivideVectors(SimpleMemory).0._State_3\);
    -- Signals:
    Signal \SimdCalculator::DivideVectors(SimpleMemory).0._Finished\: boolean := false;
    Signal \SimdCalculator::DivideVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).operation.parameter.Out.0\: \Hast.Samples.SampleAssembly.SimdOperation\;
    Signal \SimdCalculator::DivideVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\: boolean := false;
    Signal \SimdCalculator::DivideVectors(SimpleMemory).0._Started\: boolean := false;
    Signal \SimdCalculator::DivideVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\: boolean := false;
    -- System.Void Hast.Samples.SampleAssembly.SimdCalculator::DivideVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations end


    -- System.Void Hast.Samples.SampleAssembly.SimdCalculator::RunSimdOperation(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,Hast.Samples.SampleAssembly.SimdOperation).0 declarations start
    -- State machine states:
    type \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._States\ is (
        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_0\, 
        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_1\, 
        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_2\, 
        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_3\, 
        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_4\, 
        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_5\, 
        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_6\, 
        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_7\, 
        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_8\, 
        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_9\, 
        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_10\, 
        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_11\, 
        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_12\, 
        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_13\, 
        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_14\, 
        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_15\, 
        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_16\, 
        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_17\, 
        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_18\, 
        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_19\);
    -- Signals:
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._Finished\: boolean := false;
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.ReadEnable\: boolean := false;
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.WriteEnable\: boolean := false;
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.13\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.14\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.15\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.16\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.17\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.18\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.19\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.20\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.21\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.22\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.23\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.24\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.25\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.26\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.27\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.28\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.29\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.30\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.31\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.32\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.33\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.34\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.35\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.36\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.37\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.38\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.39\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.40\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.41\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.42\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.43\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.44\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.45\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.46\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.47\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.48\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.49\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.50\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.51\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.52\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.53\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.54\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.55\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.56\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.57\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.58\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.59\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.60\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.61\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.62\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.63\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.64\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.65\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.66\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.67\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.68\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.69\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.70\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.71\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.72\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.73\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.74\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.75\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.76\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.77\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.78\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.79\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.80\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.81\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.82\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.83\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.84\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.85\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.86\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.87\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.88\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.89\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.90\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.91\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.92\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.93\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.94\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.95\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.96\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.97\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.98\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.99\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.100\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.101\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.102\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.103\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.104\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.105\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.106\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.107\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.108\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.109\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.110\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.111\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.112\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.113\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.114\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.115\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.116\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.117\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.118\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.119\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.120\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.121\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.122\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.123\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.124\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.125\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.126\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.127\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.128\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.129\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.130\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.131\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.132\: signed(31 downto 0) := to_signed(0, 32);
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._Started\: boolean := false;
    Signal \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.operation.parameter.In\: \Hast.Samples.SampleAssembly.SimdOperation\;
    -- System.Void Hast.Samples.SampleAssembly.SimdCalculator::RunSimdOperation(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,Hast.Samples.SampleAssembly.SimdOperation).0 declarations end


    -- System.Void Hast::ExternalInvocationProxy() declarations start
    -- Signals:
    Signal \FinishedInternal\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ParallelAlgorithm::Run(SimpleMemory)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ObjectOrientedShowcase::Run(SimpleMemory)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumberAsync(SimpleMemory)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().PrimeCalculator::ArePrimeNumbers(SimpleMemory)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().RecursiveAlgorithms::CalculateFactorial(SimpleMemory)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().SimdCalculator::AddVectors(SimpleMemory)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().SimdCalculator::SubtractVectors(SimpleMemory)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().SimdCalculator::MultiplyVectors(SimpleMemory)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().SimdCalculator::DivideVectors(SimpleMemory)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ParallelAlgorithm::Run(SimpleMemory)._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ObjectOrientedShowcase::Run(SimpleMemory)._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumberAsync(SimpleMemory)._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().PrimeCalculator::ArePrimeNumbers(SimpleMemory)._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory)._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory)._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().RecursiveAlgorithms::CalculateFactorial(SimpleMemory)._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().SimdCalculator::AddVectors(SimpleMemory)._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().SimdCalculator::SubtractVectors(SimpleMemory)._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().SimdCalculator::MultiplyVectors(SimpleMemory)._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().SimdCalculator::DivideVectors(SimpleMemory)._Finished.0\: boolean := false;
    -- System.Void Hast::ExternalInvocationProxy() declarations end


    -- \System.Void Hast::InternalInvocationProxy()._CommonDeclarations\ declarations start
    type \InternalInvocationProxy_boolean_Array\ is array (integer range <>) of boolean;
    type \Hast::InternalInvocationProxy()._RunningStates\ is (
        WaitingForStarted, 
        WaitingForFinished, 
        AfterFinished);
    -- \System.Void Hast::InternalInvocationProxy()._CommonDeclarations\ declarations end

begin 

    -- System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32).0 state machine start
    \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._StateMachine\: process (\Clock\) 
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State\: \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._States\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_0\;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.indexObject\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.num2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.flag\: boolean := false;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.i\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.flag2\: boolean := false;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.2\: boolean := false;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.3\: boolean := false;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.4\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.5\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.6\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._Finished\ <= false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.return\ <= to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_0\;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.indexObject\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.num\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.num2\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.flag\ := false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.i\ := to_signed(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.flag2\ := false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.0\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.1\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.2\ := false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.3\ := false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.4\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.5\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.6\ := to_signed(0, 32);
            else 
                case \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State\ is 
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._Started\ = true) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._Started\ = true) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._Finished\ <= true;
                        else 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._Finished\ <= false;
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_2\ => 
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.indexObject\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.indexObject.parameter.In\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.num\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.indexObject\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.0\ := resize(\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.num\ * to_unsigned(2, 32), 32);
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.1\ := \System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::input\ + \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.0\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.num2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.1\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.flag\ := True;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.i\ := to_signed(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.i\ < to_signed(9999999, 32);
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.2\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_3\;
                        else 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_3\ => 
                        -- Repeated state of the while loop which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_2\.
                        -- The while loop's condition:
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.3\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.i\ < to_signed(9999999, 32);
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.3\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.flag2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.flag\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_6\ and ends in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_6\.
                            --     * The false branch starts in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_7\ and ends in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_7\.
                            --     * Execution after either branch will continue in the following state: \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_5\.

                            if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.flag2\) then 
                                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_6\;
                            else 
                                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_7\;
                            end if;
                        else 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_4\ => 
                        -- State after the while loop which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_2\.
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.return\ <= \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.num2\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_5\ => 
                        -- State after the if-else which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_3\.
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.flag\ := not(\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.flag\);
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.6\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.i\ + to_signed(1, 32);
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.i\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.6\;
                        -- Returning to the repeated state of the while loop which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_2\ if the loop wasn't exited with a state change.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State\ = \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_5\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_6\ => 
                        -- True branch of the if-else started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_3\.
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.4\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.num2\ + \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.num\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.num2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.4\;
                        -- Going to the state after the if-else which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_3\.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State\ = \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_6\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_7\ => 
                        -- False branch of the if-else started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_3\.
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.5\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.num2\ - \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.num\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.num2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.binaryOperationResult.5\;
                        -- Going to the state after the if-else which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_3\.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State\ = \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_7\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32).0 state machine end


    -- System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32).1 state machine start
    \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._StateMachine\: process (\Clock\) 
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State\: \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._States\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_0\;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.indexObject\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.num2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.flag\: boolean := false;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.i\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.flag2\: boolean := false;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.2\: boolean := false;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.3\: boolean := false;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.4\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.5\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.6\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._Finished\ <= false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.return\ <= to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_0\;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.indexObject\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.num\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.num2\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.flag\ := false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.i\ := to_signed(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.flag2\ := false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.0\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.1\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.2\ := false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.3\ := false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.4\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.5\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.6\ := to_signed(0, 32);
            else 
                case \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State\ is 
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._Started\ = true) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._Started\ = true) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._Finished\ <= true;
                        else 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._Finished\ <= false;
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_2\ => 
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.indexObject\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.indexObject.parameter.In\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.num\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.indexObject\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.0\ := resize(\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.num\ * to_unsigned(2, 32), 32);
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.1\ := \System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::input\ + \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.0\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.num2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.1\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.flag\ := True;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.i\ := to_signed(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.i\ < to_signed(9999999, 32);
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.2\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_3\;
                        else 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_3\ => 
                        -- Repeated state of the while loop which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_2\.
                        -- The while loop's condition:
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.3\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.i\ < to_signed(9999999, 32);
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.3\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.flag2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.flag\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_6\ and ends in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_6\.
                            --     * The false branch starts in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_7\ and ends in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_7\.
                            --     * Execution after either branch will continue in the following state: \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_5\.

                            if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.flag2\) then 
                                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_6\;
                            else 
                                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_7\;
                            end if;
                        else 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_4\ => 
                        -- State after the while loop which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_2\.
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.return\ <= \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.num2\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_5\ => 
                        -- State after the if-else which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_3\.
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.flag\ := not(\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.flag\);
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.6\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.i\ + to_signed(1, 32);
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.i\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.6\;
                        -- Returning to the repeated state of the while loop which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_2\ if the loop wasn't exited with a state change.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State\ = \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_5\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_6\ => 
                        -- True branch of the if-else started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_3\.
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.4\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.num2\ + \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.num\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.num2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.4\;
                        -- Going to the state after the if-else which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_3\.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State\ = \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_6\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_7\ => 
                        -- False branch of the if-else started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_3\.
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.5\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.num2\ - \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.num\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.num2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.binaryOperationResult.5\;
                        -- Going to the state after the if-else which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_3\.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State\ = \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_7\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32).1 state machine end


    -- System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32).2 state machine start
    \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._StateMachine\: process (\Clock\) 
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State\: \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._States\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_0\;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.indexObject\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.num2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.flag\: boolean := false;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.i\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.flag2\: boolean := false;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.2\: boolean := false;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.3\: boolean := false;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.4\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.5\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.6\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._Finished\ <= false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.return\ <= to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_0\;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.indexObject\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.num\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.num2\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.flag\ := false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.i\ := to_signed(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.flag2\ := false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.0\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.1\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.2\ := false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.3\ := false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.4\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.5\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.6\ := to_signed(0, 32);
            else 
                case \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State\ is 
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._Started\ = true) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._Started\ = true) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._Finished\ <= true;
                        else 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._Finished\ <= false;
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_2\ => 
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.indexObject\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.indexObject.parameter.In\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.num\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.indexObject\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.0\ := resize(\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.num\ * to_unsigned(2, 32), 32);
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.1\ := \System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::input\ + \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.0\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.num2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.1\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.flag\ := True;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.i\ := to_signed(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.i\ < to_signed(9999999, 32);
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.2\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_3\;
                        else 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_3\ => 
                        -- Repeated state of the while loop which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_2\.
                        -- The while loop's condition:
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.3\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.i\ < to_signed(9999999, 32);
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.3\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.flag2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.flag\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_6\ and ends in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_6\.
                            --     * The false branch starts in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_7\ and ends in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_7\.
                            --     * Execution after either branch will continue in the following state: \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_5\.

                            if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.flag2\) then 
                                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_6\;
                            else 
                                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_7\;
                            end if;
                        else 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_4\ => 
                        -- State after the while loop which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_2\.
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.return\ <= \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.num2\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_5\ => 
                        -- State after the if-else which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_3\.
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.flag\ := not(\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.flag\);
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.6\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.i\ + to_signed(1, 32);
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.i\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.6\;
                        -- Returning to the repeated state of the while loop which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_2\ if the loop wasn't exited with a state change.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State\ = \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_5\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_6\ => 
                        -- True branch of the if-else started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_3\.
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.4\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.num2\ + \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.num\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.num2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.4\;
                        -- Going to the state after the if-else which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_3\.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State\ = \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_6\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_7\ => 
                        -- False branch of the if-else started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_3\.
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.5\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.num2\ - \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.num\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.num2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.binaryOperationResult.5\;
                        -- Going to the state after the if-else which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_3\.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State\ = \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_7\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32).2 state machine end


    -- System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32).3 state machine start
    \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._StateMachine\: process (\Clock\) 
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State\: \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._States\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_0\;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.indexObject\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.num2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.flag\: boolean := false;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.i\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.flag2\: boolean := false;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.2\: boolean := false;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.3\: boolean := false;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.4\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.5\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.6\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._Finished\ <= false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.return\ <= to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_0\;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.indexObject\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.num\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.num2\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.flag\ := false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.i\ := to_signed(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.flag2\ := false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.0\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.1\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.2\ := false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.3\ := false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.4\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.5\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.6\ := to_signed(0, 32);
            else 
                case \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State\ is 
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._Started\ = true) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._Started\ = true) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._Finished\ <= true;
                        else 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._Finished\ <= false;
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_2\ => 
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.indexObject\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.indexObject.parameter.In\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.num\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.indexObject\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.0\ := resize(\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.num\ * to_unsigned(2, 32), 32);
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.1\ := \System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::input\ + \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.0\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.num2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.1\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.flag\ := True;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.i\ := to_signed(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.i\ < to_signed(9999999, 32);
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.2\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_3\;
                        else 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_3\ => 
                        -- Repeated state of the while loop which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_2\.
                        -- The while loop's condition:
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.3\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.i\ < to_signed(9999999, 32);
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.3\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.flag2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.flag\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_6\ and ends in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_6\.
                            --     * The false branch starts in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_7\ and ends in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_7\.
                            --     * Execution after either branch will continue in the following state: \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_5\.

                            if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.flag2\) then 
                                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_6\;
                            else 
                                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_7\;
                            end if;
                        else 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_4\ => 
                        -- State after the while loop which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_2\.
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.return\ <= \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.num2\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_5\ => 
                        -- State after the if-else which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_3\.
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.flag\ := not(\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.flag\);
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.6\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.i\ + to_signed(1, 32);
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.i\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.6\;
                        -- Returning to the repeated state of the while loop which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_2\ if the loop wasn't exited with a state change.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State\ = \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_5\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_6\ => 
                        -- True branch of the if-else started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_3\.
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.4\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.num2\ + \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.num\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.num2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.4\;
                        -- Going to the state after the if-else which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_3\.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State\ = \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_6\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_7\ => 
                        -- False branch of the if-else started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_3\.
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.5\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.num2\ - \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.num\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.num2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.binaryOperationResult.5\;
                        -- Going to the state after the if-else which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_3\.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State\ = \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_7\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32).3 state machine end


    -- System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32).4 state machine start
    \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._StateMachine\: process (\Clock\) 
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State\: \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._States\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_0\;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.indexObject\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.num2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.flag\: boolean := false;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.i\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.flag2\: boolean := false;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.2\: boolean := false;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.3\: boolean := false;
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.4\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.5\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.6\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._Finished\ <= false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.return\ <= to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_0\;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.indexObject\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.num\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.num2\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.flag\ := false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.i\ := to_signed(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.flag2\ := false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.0\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.1\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.2\ := false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.3\ := false;
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.4\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.5\ := to_unsigned(0, 32);
                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.6\ := to_signed(0, 32);
            else 
                case \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State\ is 
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._Started\ = true) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._Started\ = true) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._Finished\ <= true;
                        else 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._Finished\ <= false;
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_2\ => 
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.indexObject\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.indexObject.parameter.In\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.num\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.indexObject\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.0\ := resize(\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.num\ * to_unsigned(2, 32), 32);
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.1\ := \System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::input\ + \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.0\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.num2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.1\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.flag\ := True;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.i\ := to_signed(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.i\ < to_signed(9999999, 32);
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.2\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_3\;
                        else 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_3\ => 
                        -- Repeated state of the while loop which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_2\.
                        -- The while loop's condition:
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.3\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.i\ < to_signed(9999999, 32);
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.3\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.flag2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.flag\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_6\ and ends in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_6\.
                            --     * The false branch starts in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_7\ and ends in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_7\.
                            --     * Execution after either branch will continue in the following state: \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_5\.

                            if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.flag2\) then 
                                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_6\;
                            else 
                                \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_7\;
                            end if;
                        else 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_4\ => 
                        -- State after the while loop which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_2\.
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.return\ <= \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.num2\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_5\ => 
                        -- State after the if-else which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_3\.
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.flag\ := not(\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.flag\);
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.6\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.i\ + to_signed(1, 32);
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.i\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.6\;
                        -- Returning to the repeated state of the while loop which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_2\ if the loop wasn't exited with a state change.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State\ = \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_5\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_6\ => 
                        -- True branch of the if-else started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_3\.
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.4\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.num2\ + \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.num\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.num2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.4\;
                        -- Going to the state after the if-else which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_3\.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State\ = \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_6\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_7\ => 
                        -- False branch of the if-else started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_3\.
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.5\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.num2\ - \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.num\;
                        \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.num2\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.binaryOperationResult.5\;
                        -- Going to the state after the if-else which was started in state \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_3\.
                        if (\ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State\ = \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_7\) then 
                            \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State\ := \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32).4 state machine end


    -- System.Void Hast.Samples.SampleAssembly.ParallelAlgorithm::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine start
    \ParallelAlgorithm::Run(SimpleMemory).0._StateMachine\: process (\Clock\) 
        Variable \ParallelAlgorithm::Run(SimpleMemory).0._State\: \ParallelAlgorithm::Run(SimpleMemory).0._States\ := \ParallelAlgorithm::Run(SimpleMemory).0._State_0\;
        Variable \ParallelAlgorithm::Run(SimpleMemory).0.array\: \unsigned32_Array\(0 to 279) := (others => to_unsigned(0, 32));
        Variable \ParallelAlgorithm::Run(SimpleMemory).0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm::Run(SimpleMemory).0.arg_57_1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ParallelAlgorithm::Run(SimpleMemory).0.num2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm::Run(SimpleMemory).0.i\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ParallelAlgorithm::Run(SimpleMemory).0.dataIn.0\: std_logic_vector(31 downto 0);
        Variable \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.0\: boolean := false;
        Variable \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.1\: boolean := false;
        Variable \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).invocationIndex\: integer range 0 to 4 := 0;
        Variable \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm::Run(SimpleMemory).0.return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm::Run(SimpleMemory).0.return.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm::Run(SimpleMemory).0.return.2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm::Run(SimpleMemory).0.return.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm::Run(SimpleMemory).0.return.4\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.3\: boolean := false;
        Variable \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.4\: boolean := false;
        Variable \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.5\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.6\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ParallelAlgorithm::Run(SimpleMemory).0._Finished\ <= false;
                \ParallelAlgorithm::Run(SimpleMemory).0.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \ParallelAlgorithm::Run(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                \ParallelAlgorithm::Run(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).indexObject.parameter.Out.0\ <= to_unsigned(0, 32);
                \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.0\ <= false;
                \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).indexObject.parameter.Out.1\ <= to_unsigned(0, 32);
                \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.1\ <= false;
                \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).indexObject.parameter.Out.2\ <= to_unsigned(0, 32);
                \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.2\ <= false;
                \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).indexObject.parameter.Out.3\ <= to_unsigned(0, 32);
                \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.3\ <= false;
                \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).indexObject.parameter.Out.4\ <= to_unsigned(0, 32);
                \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.4\ <= false;
                \ParallelAlgorithm::Run(SimpleMemory).0._State\ := \ParallelAlgorithm::Run(SimpleMemory).0._State_0\;
                \ParallelAlgorithm::Run(SimpleMemory).0.array\ := (others => to_unsigned(0, 32));
                \ParallelAlgorithm::Run(SimpleMemory).0.num\ := to_unsigned(0, 32);
                \ParallelAlgorithm::Run(SimpleMemory).0.arg_57_1\ := to_signed(0, 32);
                \ParallelAlgorithm::Run(SimpleMemory).0.num2\ := to_unsigned(0, 32);
                \ParallelAlgorithm::Run(SimpleMemory).0.i\ := to_signed(0, 32);
                \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.0\ := false;
                \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.1\ := false;
                \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).invocationIndex\ := 0;
                \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.2\ := to_unsigned(0, 32);
                \ParallelAlgorithm::Run(SimpleMemory).0.return.0\ := to_unsigned(0, 32);
                \ParallelAlgorithm::Run(SimpleMemory).0.return.1\ := to_unsigned(0, 32);
                \ParallelAlgorithm::Run(SimpleMemory).0.return.2\ := to_unsigned(0, 32);
                \ParallelAlgorithm::Run(SimpleMemory).0.return.3\ := to_unsigned(0, 32);
                \ParallelAlgorithm::Run(SimpleMemory).0.return.4\ := to_unsigned(0, 32);
                \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.3\ := false;
                \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.4\ := false;
                \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.5\ := to_unsigned(0, 32);
                \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.6\ := to_signed(0, 32);
            else 
                case \ParallelAlgorithm::Run(SimpleMemory).0._State\ is 
                    when \ParallelAlgorithm::Run(SimpleMemory).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ParallelAlgorithm::Run(SimpleMemory).0._Started\ = true) then 
                            \ParallelAlgorithm::Run(SimpleMemory).0._State\ := \ParallelAlgorithm::Run(SimpleMemory).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelAlgorithm::Run(SimpleMemory).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ParallelAlgorithm::Run(SimpleMemory).0._Started\ = true) then 
                            \ParallelAlgorithm::Run(SimpleMemory).0._Finished\ <= true;
                        else 
                            \ParallelAlgorithm::Run(SimpleMemory).0._Finished\ <= false;
                            \ParallelAlgorithm::Run(SimpleMemory).0._State\ := \ParallelAlgorithm::Run(SimpleMemory).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelAlgorithm::Run(SimpleMemory).0._State_2\ => 
                        -- Begin SimpleMemory read.
                        \ParallelAlgorithm::Run(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(to_signed(0, 32), 32);
                        \ParallelAlgorithm::Run(SimpleMemory).0.SimpleMemory.ReadEnable\ <= true;
                        \ParallelAlgorithm::Run(SimpleMemory).0._State\ := \ParallelAlgorithm::Run(SimpleMemory).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelAlgorithm::Run(SimpleMemory).0._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \ParallelAlgorithm::Run(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                            \ParallelAlgorithm::Run(SimpleMemory).0.dataIn.0\ := \DataIn\;
                            \System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::input\ := ConvertStdLogicVectorToUInt32(\ParallelAlgorithm::Run(SimpleMemory).0.dataIn.0\);
                            \ParallelAlgorithm::Run(SimpleMemory).0.array\ := (others => to_unsigned(0, 32));
                            \ParallelAlgorithm::Run(SimpleMemory).0.num\ := to_unsigned(0, 32);
                            -- Starting a while loop.
                            -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                            \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.0\ := \ParallelAlgorithm::Run(SimpleMemory).0.num\ < to_unsigned(280, 32);
                            if (\ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.0\) then 
                                \ParallelAlgorithm::Run(SimpleMemory).0._State\ := \ParallelAlgorithm::Run(SimpleMemory).0._State_4\;
                            else 
                                \ParallelAlgorithm::Run(SimpleMemory).0._State\ := \ParallelAlgorithm::Run(SimpleMemory).0._State_5\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ParallelAlgorithm::Run(SimpleMemory).0._State_4\ => 
                        -- Repeated state of the while loop which was started in state \ParallelAlgorithm::Run(SimpleMemory).0._State_3\.
                        -- The while loop's condition:
                        \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.1\ := \ParallelAlgorithm::Run(SimpleMemory).0.num\ < to_unsigned(280, 32);
                        if (\ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.1\) then 
                            \ParallelAlgorithm::Run(SimpleMemory).0.arg_57_1\ := signed(\ParallelAlgorithm::Run(SimpleMemory).0.num\);
                            -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32)
                            case \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).invocationIndex\ is 
                                when 0 => 
                                    \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).indexObject.parameter.Out.0\ <= \ParallelAlgorithm::Run(SimpleMemory).0.num\;
                                    \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.0\ <= true;
                                when 1 => 
                                    \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).indexObject.parameter.Out.1\ <= \ParallelAlgorithm::Run(SimpleMemory).0.num\;
                                    \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.1\ <= true;
                                when 2 => 
                                    \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).indexObject.parameter.Out.2\ <= \ParallelAlgorithm::Run(SimpleMemory).0.num\;
                                    \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.2\ <= true;
                                when 3 => 
                                    \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).indexObject.parameter.Out.3\ <= \ParallelAlgorithm::Run(SimpleMemory).0.num\;
                                    \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.3\ <= true;
                                when 4 => 
                                    \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).indexObject.parameter.Out.4\ <= \ParallelAlgorithm::Run(SimpleMemory).0.num\;
                                    \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.4\ <= true;
                            end case;
                            \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).invocationIndex\ := \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).invocationIndex\ + 1;
                            \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.2\ := \ParallelAlgorithm::Run(SimpleMemory).0.num\ + to_unsigned(1, 32);
                            \ParallelAlgorithm::Run(SimpleMemory).0.num\ := \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.2\;
                        else 
                            \ParallelAlgorithm::Run(SimpleMemory).0._State\ := \ParallelAlgorithm::Run(SimpleMemory).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \ParallelAlgorithm::Run(SimpleMemory).0._State_5\ => 
                        -- State after the while loop which was started in state \ParallelAlgorithm::Run(SimpleMemory).0._State_3\.
                        \ParallelAlgorithm::Run(SimpleMemory).0._State\ := \ParallelAlgorithm::Run(SimpleMemory).0._State_6\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelAlgorithm::Run(SimpleMemory).0._State_6\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32)
                        if (\ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.1\ = \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Finished.1\ and \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.2\ = \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Finished.2\ and \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.3\ = \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Finished.3\ and \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.4\ = \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Finished.4\ and \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.0\ = \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Finished.0\) then 
                            \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.0\ <= false;
                            \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.1\ <= false;
                            \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.2\ <= false;
                            \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.3\ <= false;
                            \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.4\ <= false;
                            \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).invocationIndex\ := 0;
                            \ParallelAlgorithm::Run(SimpleMemory).0.return.0\ := \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).return.0\;
                            \ParallelAlgorithm::Run(SimpleMemory).0.return.1\ := \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).return.1\;
                            \ParallelAlgorithm::Run(SimpleMemory).0.return.2\ := \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).return.2\;
                            \ParallelAlgorithm::Run(SimpleMemory).0.return.3\ := \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).return.3\;
                            \ParallelAlgorithm::Run(SimpleMemory).0.return.4\ := \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).return.4\;
                            \ParallelAlgorithm::Run(SimpleMemory).0.array\(0) := \ParallelAlgorithm::Run(SimpleMemory).0.return.0\;
                            \ParallelAlgorithm::Run(SimpleMemory).0.array\(1) := \ParallelAlgorithm::Run(SimpleMemory).0.return.1\;
                            \ParallelAlgorithm::Run(SimpleMemory).0.array\(2) := \ParallelAlgorithm::Run(SimpleMemory).0.return.2\;
                            \ParallelAlgorithm::Run(SimpleMemory).0.array\(3) := \ParallelAlgorithm::Run(SimpleMemory).0.return.3\;
                            \ParallelAlgorithm::Run(SimpleMemory).0.array\(4) := \ParallelAlgorithm::Run(SimpleMemory).0.return.4\;
                            \ParallelAlgorithm::Run(SimpleMemory).0.num2\ := to_unsigned(0, 32);
                            \ParallelAlgorithm::Run(SimpleMemory).0.i\ := to_signed(0, 32);
                            -- Starting a while loop.
                            -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                            \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.3\ := \ParallelAlgorithm::Run(SimpleMemory).0.i\ < to_signed(280, 32);
                            if (\ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.3\) then 
                                \ParallelAlgorithm::Run(SimpleMemory).0._State\ := \ParallelAlgorithm::Run(SimpleMemory).0._State_7\;
                            else 
                                \ParallelAlgorithm::Run(SimpleMemory).0._State\ := \ParallelAlgorithm::Run(SimpleMemory).0._State_8\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ParallelAlgorithm::Run(SimpleMemory).0._State_7\ => 
                        -- Repeated state of the while loop which was started in state \ParallelAlgorithm::Run(SimpleMemory).0._State_6\.
                        -- The while loop's condition:
                        \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.4\ := \ParallelAlgorithm::Run(SimpleMemory).0.i\ < to_signed(280, 32);
                        if (\ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.4\) then 
                            \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.5\ := \ParallelAlgorithm::Run(SimpleMemory).0.num2\ + \ParallelAlgorithm::Run(SimpleMemory).0.array\(to_integer(\ParallelAlgorithm::Run(SimpleMemory).0.i\));
                            \ParallelAlgorithm::Run(SimpleMemory).0.num2\ := \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.5\;
                            \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.6\ := \ParallelAlgorithm::Run(SimpleMemory).0.i\ + to_signed(1, 32);
                            \ParallelAlgorithm::Run(SimpleMemory).0.i\ := \ParallelAlgorithm::Run(SimpleMemory).0.binaryOperationResult.6\;
                        else 
                            \ParallelAlgorithm::Run(SimpleMemory).0._State\ := \ParallelAlgorithm::Run(SimpleMemory).0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \ParallelAlgorithm::Run(SimpleMemory).0._State_8\ => 
                        -- State after the while loop which was started in state \ParallelAlgorithm::Run(SimpleMemory).0._State_6\.
                        -- Begin SimpleMemory write.
                        \ParallelAlgorithm::Run(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(to_signed(0, 32), 32);
                        \ParallelAlgorithm::Run(SimpleMemory).0.SimpleMemory.WriteEnable\ <= true;
                        \ParallelAlgorithm::Run(SimpleMemory).0.SimpleMemory.DataOut\ <= ConvertUInt32ToStdLogicVector(\ParallelAlgorithm::Run(SimpleMemory).0.num2\);
                        \ParallelAlgorithm::Run(SimpleMemory).0._State\ := \ParallelAlgorithm::Run(SimpleMemory).0._State_9\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelAlgorithm::Run(SimpleMemory).0._State_9\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \ParallelAlgorithm::Run(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                            \ParallelAlgorithm::Run(SimpleMemory).0._State\ := \ParallelAlgorithm::Run(SimpleMemory).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.Samples.SampleAssembly.ParallelAlgorithm::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine end


    -- System.Void Hast.Samples.SampleAssembly.ObjectOrientedShowcase::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine start
    \ObjectOrientedShowcase::Run(SimpleMemory).0._StateMachine\: process (\Clock\) 
        Variable \ObjectOrientedShowcase::Run(SimpleMemory).0._State\: \ObjectOrientedShowcase::Run(SimpleMemory).0._States\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_0\;
        Variable \ObjectOrientedShowcase::Run(SimpleMemory).0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ObjectOrientedShowcase::Run(SimpleMemory).0.array\: \Hast.Samples.SampleAssembly.NumberContainer_Array\(0 to 3);
        Variable \ObjectOrientedShowcase::Run(SimpleMemory).0.array2\: \Hast.Samples.SampleAssembly.NumberContainer_Array\(0 to 0);
        Variable \ObjectOrientedShowcase::Run(SimpleMemory).0.numberContainer\: \Hast.Samples.SampleAssembly.NumberContainer\;
        Variable \ObjectOrientedShowcase::Run(SimpleMemory).0.flag\: boolean := false;
        Variable \ObjectOrientedShowcase::Run(SimpleMemory).0.i\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ObjectOrientedShowcase::Run(SimpleMemory).0.dataIn.0\: std_logic_vector(31 downto 0);
        Variable \ObjectOrientedShowcase::Run(SimpleMemory).0.object29a6fc5705986afeb93844c5d0476ea3403f870b46cc8be7ca071f85ea3d7508\: \Hast.Samples.SampleAssembly.MemoryContainer\;
        Variable \ObjectOrientedShowcase::Run(SimpleMemory).0.return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ObjectOrientedShowcase::Run(SimpleMemory).0.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ObjectOrientedShowcase::Run(SimpleMemory).0.binaryOperationResult.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ObjectOrientedShowcase::Run(SimpleMemory).0.return.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ObjectOrientedShowcase::Run(SimpleMemory).0.return.2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ObjectOrientedShowcase::Run(SimpleMemory).0.return.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ObjectOrientedShowcase::Run(SimpleMemory).0.binaryOperationResult.2\: boolean := false;
        Variable \ObjectOrientedShowcase::Run(SimpleMemory).0.binaryOperationResult.3\: boolean := false;
        Variable \ObjectOrientedShowcase::Run(SimpleMemory).0.return.4\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ObjectOrientedShowcase::Run(SimpleMemory).0.binaryOperationResult.4\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ObjectOrientedShowcase::Run(SimpleMemory).0.return.5\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ObjectOrientedShowcase::Run(SimpleMemory).0._Finished\ <= false;
                \ObjectOrientedShowcase::Run(SimpleMemory).0.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \ObjectOrientedShowcase::Run(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                \ObjectOrientedShowcase::Run(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::.ctor(SimpleMemory)._Started.0\ <= false;
                \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::GetInput()._Started.0\ <= false;
                \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor()._Started.0\ <= false;
                \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor(UInt32).number.parameter.Out.0\ <= to_unsigned(0, 32);
                \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor(UInt32)._Started.0\ <= false;
                \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::set_NumberPlusFive(UInt32).value.parameter.Out.0\ <= to_unsigned(0, 32);
                \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::set_NumberPlusFive(UInt32)._Started.0\ <= false;
                \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32).increaseBy.parameter.Out.0\ <= to_unsigned(0, 32);
                \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32)._Started.0\ <= false;
                \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::get_NumberPlusFive()._Started.0\ <= false;
                \ObjectOrientedShowcase::Run(SimpleMemory).0.ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[])._Started.0\ <= false;
                \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_0\;
                \ObjectOrientedShowcase::Run(SimpleMemory).0.num\ := to_unsigned(0, 32);
                \ObjectOrientedShowcase::Run(SimpleMemory).0.flag\ := false;
                \ObjectOrientedShowcase::Run(SimpleMemory).0.i\ := to_signed(0, 32);
                \ObjectOrientedShowcase::Run(SimpleMemory).0.return.0\ := to_unsigned(0, 32);
                \ObjectOrientedShowcase::Run(SimpleMemory).0.binaryOperationResult.0\ := to_unsigned(0, 32);
                \ObjectOrientedShowcase::Run(SimpleMemory).0.binaryOperationResult.1\ := to_unsigned(0, 32);
                \ObjectOrientedShowcase::Run(SimpleMemory).0.return.1\ := to_unsigned(0, 32);
                \ObjectOrientedShowcase::Run(SimpleMemory).0.return.2\ := to_unsigned(0, 32);
                \ObjectOrientedShowcase::Run(SimpleMemory).0.return.3\ := to_unsigned(0, 32);
                \ObjectOrientedShowcase::Run(SimpleMemory).0.binaryOperationResult.2\ := false;
                \ObjectOrientedShowcase::Run(SimpleMemory).0.binaryOperationResult.3\ := false;
                \ObjectOrientedShowcase::Run(SimpleMemory).0.return.4\ := to_unsigned(0, 32);
                \ObjectOrientedShowcase::Run(SimpleMemory).0.binaryOperationResult.4\ := to_signed(0, 32);
                \ObjectOrientedShowcase::Run(SimpleMemory).0.return.5\ := to_unsigned(0, 32);
            else 
                case \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ is 
                    when \ObjectOrientedShowcase::Run(SimpleMemory).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ObjectOrientedShowcase::Run(SimpleMemory).0._Started\ = true) then 
                            \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectOrientedShowcase::Run(SimpleMemory).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ObjectOrientedShowcase::Run(SimpleMemory).0._Started\ = true) then 
                            \ObjectOrientedShowcase::Run(SimpleMemory).0._Finished\ <= true;
                        else 
                            \ObjectOrientedShowcase::Run(SimpleMemory).0._Finished\ <= false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectOrientedShowcase::Run(SimpleMemory).0._State_2\ => 
                        -- Begin SimpleMemory read.
                        \ObjectOrientedShowcase::Run(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(to_signed(0, 32), 32);
                        \ObjectOrientedShowcase::Run(SimpleMemory).0.SimpleMemory.ReadEnable\ <= true;
                        \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectOrientedShowcase::Run(SimpleMemory).0._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.dataIn.0\ := \DataIn\;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.num\ := ConvertStdLogicVectorToUInt32(\ObjectOrientedShowcase::Run(SimpleMemory).0.dataIn.0\);
                            -- Initializing record fields to their defaults.
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.object29a6fc5705986afeb93844c5d0476ea3403f870b46cc8be7ca071f85ea3d7508\.\IsNull\ := false;
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Hast.Samples.SampleAssembly.MemoryContainer::.ctor(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory)
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::.ctor(SimpleMemory).this.parameter.Out.0\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.object29a6fc5705986afeb93844c5d0476ea3403f870b46cc8be7ca071f85ea3d7508\;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::.ctor(SimpleMemory)._Started.0\ <= true;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectOrientedShowcase::Run(SimpleMemory).0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.Samples.SampleAssembly.MemoryContainer::.ctor(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory)
                        if (\ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::.ctor(SimpleMemory)._Started.0\ = \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::.ctor(SimpleMemory)._Finished.0\) then 
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::.ctor(SimpleMemory)._Started.0\ <= false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.object29a6fc5705986afeb93844c5d0476ea3403f870b46cc8be7ca071f85ea3d7508\ := \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::.ctor(SimpleMemory).this.parameter.In.0\;
                            -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.MemoryContainer::GetInput()
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::GetInput().this.parameter.Out.0\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.object29a6fc5705986afeb93844c5d0476ea3403f870b46cc8be7ca071f85ea3d7508\;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::GetInput()._Started.0\ <= true;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectOrientedShowcase::Run(SimpleMemory).0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.MemoryContainer::GetInput()
                        if (\ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::GetInput()._Started.0\ = \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::GetInput()._Finished.0\) then 
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::GetInput()._Started.0\ <= false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.return.0\ := \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::GetInput().return.0\;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.object29a6fc5705986afeb93844c5d0476ea3403f870b46cc8be7ca071f85ea3d7508\ := \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::GetInput().this.parameter.In.0\;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.num\ := \ObjectOrientedShowcase::Run(SimpleMemory).0.return.0\;
                            -- Initializing record fields to their defaults.
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(0, 32))).\IsNull\ := false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(0, 32))).\WasIncreased\ := false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(0, 32))).\Number\ := to_unsigned(0, 32);
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Hast.Samples.SampleAssembly.NumberContainer::.ctor()
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor().this.parameter.Out.0\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(0, 32)));
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor()._Started.0\ <= true;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectOrientedShowcase::Run(SimpleMemory).0._State_6\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.Samples.SampleAssembly.NumberContainer::.ctor()
                        if (\ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor()._Started.0\ = \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor()._Finished.0\) then 
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor()._Started.0\ <= false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(0, 32))) := \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor().this.parameter.In.0\;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(0, 32))).\Number\ := \ObjectOrientedShowcase::Run(SimpleMemory).0.num\;
                            -- Initializing record fields to their defaults.
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(1, 32))).\IsNull\ := false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(1, 32))).\WasIncreased\ := false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(1, 32))).\Number\ := to_unsigned(0, 32);
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Hast.Samples.SampleAssembly.NumberContainer::.ctor()
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor().this.parameter.Out.0\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(1, 32)));
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor()._Started.0\ <= true;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectOrientedShowcase::Run(SimpleMemory).0._State_7\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.Samples.SampleAssembly.NumberContainer::.ctor()
                        if (\ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor()._Started.0\ = \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor()._Finished.0\) then 
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor()._Started.0\ <= false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(1, 32))) := \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor().this.parameter.In.0\;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.binaryOperationResult.0\ := \ObjectOrientedShowcase::Run(SimpleMemory).0.num\ + to_unsigned(4, 32);
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(1, 32))).\Number\ := \ObjectOrientedShowcase::Run(SimpleMemory).0.binaryOperationResult.0\;
                            -- Initializing record fields to their defaults.
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(2, 32))).\IsNull\ := false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(2, 32))).\WasIncreased\ := false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(2, 32))).\Number\ := to_unsigned(0, 32);
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Hast.Samples.SampleAssembly.NumberContainer::.ctor()
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor().this.parameter.Out.0\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(2, 32)));
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor()._Started.0\ <= true;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ObjectOrientedShowcase::Run(SimpleMemory).0._State_8\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.Samples.SampleAssembly.NumberContainer::.ctor()
                        if (\ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor()._Started.0\ = \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor()._Finished.0\) then 
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor()._Started.0\ <= false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(2, 32))) := \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor().this.parameter.In.0\;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(2, 32))).\Number\ := to_unsigned(24, 32);
                            -- Initializing record fields to their defaults.
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(3, 32))).\IsNull\ := false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(3, 32))).\WasIncreased\ := false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(3, 32))).\Number\ := to_unsigned(0, 32);
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Hast.Samples.SampleAssembly.NumberContainer::.ctor(System.UInt32)
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor(UInt32).this.parameter.Out.0\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(3, 32)));
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor(UInt32).number.parameter.Out.0\ <= to_unsigned(9, 32);
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor(UInt32)._Started.0\ <= true;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_9\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectOrientedShowcase::Run(SimpleMemory).0._State_9\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.Samples.SampleAssembly.NumberContainer::.ctor(System.UInt32)
                        if (\ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor(UInt32)._Started.0\ = \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor(UInt32)._Finished.0\) then 
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor(UInt32)._Started.0\ <= false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(3, 32))) := \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor(UInt32).this.parameter.In.0\;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.binaryOperationResult.1\ := \ObjectOrientedShowcase::Run(SimpleMemory).0.num\ + to_unsigned(10, 32);
                            -- Starting state machine invocation for the following method: System.Void Hast.Samples.SampleAssembly.NumberContainer::set_NumberPlusFive(System.UInt32)
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::set_NumberPlusFive(UInt32).this.parameter.Out.0\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(0, 32)));
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::set_NumberPlusFive(UInt32).value.parameter.Out.0\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.binaryOperationResult.1\;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::set_NumberPlusFive(UInt32)._Started.0\ <= true;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_10\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ObjectOrientedShowcase::Run(SimpleMemory).0._State_10\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.Samples.SampleAssembly.NumberContainer::set_NumberPlusFive(System.UInt32)
                        if (\ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::set_NumberPlusFive(UInt32)._Started.0\ = \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::set_NumberPlusFive(UInt32)._Finished.0\) then 
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::set_NumberPlusFive(UInt32)._Started.0\ <= false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(0, 32))) := \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::set_NumberPlusFive(UInt32).this.parameter.In.0\;
                            -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.NumberContainer::IncreaseNumber(System.UInt32)
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32).this.parameter.Out.0\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(1, 32)));
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32).increaseBy.parameter.Out.0\ <= to_unsigned(5, 32);
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32)._Started.0\ <= true;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_11\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectOrientedShowcase::Run(SimpleMemory).0._State_11\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.NumberContainer::IncreaseNumber(System.UInt32)
                        if (\ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32)._Started.0\ = \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32)._Finished.0\) then 
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32)._Started.0\ <= false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.return.1\ := \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32).return.0\;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(to_signed(1, 32))) := \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32).this.parameter.In.0\;
                            -- Initializing record fields to their defaults.
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.numberContainer\.\IsNull\ := false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.numberContainer\.\WasIncreased\ := false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.numberContainer\.\Number\ := to_unsigned(0, 32);
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Hast.Samples.SampleAssembly.NumberContainer::.ctor()
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor().this.parameter.Out.0\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.numberContainer\;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor()._Started.0\ <= true;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_12\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectOrientedShowcase::Run(SimpleMemory).0._State_12\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.Samples.SampleAssembly.NumberContainer::.ctor()
                        if (\ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor()._Started.0\ = \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor()._Finished.0\) then 
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor()._Started.0\ <= false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.numberContainer\ := \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor().this.parameter.In.0\;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.numberContainer\.\Number\ := to_unsigned(5, 32);
                            -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.NumberContainer::get_NumberPlusFive()
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::get_NumberPlusFive().this.parameter.Out.0\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.numberContainer\;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::get_NumberPlusFive()._Started.0\ <= true;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_13\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectOrientedShowcase::Run(SimpleMemory).0._State_13\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.NumberContainer::get_NumberPlusFive()
                        if (\ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::get_NumberPlusFive()._Started.0\ = \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::get_NumberPlusFive()._Finished.0\) then 
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::get_NumberPlusFive()._Started.0\ <= false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.return.2\ := \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::get_NumberPlusFive().return.0\;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.numberContainer\ := \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::get_NumberPlusFive().this.parameter.In.0\;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.numberContainer\.\Number\ := \ObjectOrientedShowcase::Run(SimpleMemory).0.return.2\;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.flag\ := not(\ObjectOrientedShowcase::Run(SimpleMemory).0.numberContainer\.\WasIncreased\);

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \ObjectOrientedShowcase::Run(SimpleMemory).0._State_15\ and ends in state \ObjectOrientedShowcase::Run(SimpleMemory).0._State_16\.
                            --     * Execution after either branch will continue in the following state: \ObjectOrientedShowcase::Run(SimpleMemory).0._State_14\.

                            if (\ObjectOrientedShowcase::Run(SimpleMemory).0.flag\) then 
                                \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_15\;
                            else 
                                -- There was no false branch, so going directly to the state after the if-else.
                                \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_14\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ObjectOrientedShowcase::Run(SimpleMemory).0._State_14\ => 
                        -- State after the if-else which was started in state \ObjectOrientedShowcase::Run(SimpleMemory).0._State_13\.
                        \ObjectOrientedShowcase::Run(SimpleMemory).0.array2\(to_integer(to_signed(0, 32))) := \ObjectOrientedShowcase::Run(SimpleMemory).0.numberContainer\;
                        \ObjectOrientedShowcase::Run(SimpleMemory).0.i\ := to_signed(0, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \ObjectOrientedShowcase::Run(SimpleMemory).0.binaryOperationResult.2\ := \ObjectOrientedShowcase::Run(SimpleMemory).0.i\ < to_signed(4, 32);
                        if (\ObjectOrientedShowcase::Run(SimpleMemory).0.binaryOperationResult.2\) then 
                            \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_17\;
                        else 
                            \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_18\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ObjectOrientedShowcase::Run(SimpleMemory).0._State_15\ => 
                        -- True branch of the if-else started in state \ObjectOrientedShowcase::Run(SimpleMemory).0._State_13\.
                        -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.NumberContainer::IncreaseNumber(System.UInt32)
                        \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32).this.parameter.Out.0\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.numberContainer\;
                        \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32).increaseBy.parameter.Out.0\ <= to_unsigned(5, 32);
                        \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32)._Started.0\ <= true;
                        \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_16\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectOrientedShowcase::Run(SimpleMemory).0._State_16\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.NumberContainer::IncreaseNumber(System.UInt32)
                        if (\ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32)._Started.0\ = \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32)._Finished.0\) then 
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32)._Started.0\ <= false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.return.3\ := \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32).return.0\;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.numberContainer\ := \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32).this.parameter.In.0\;
                            -- Going to the state after the if-else which was started in state \ObjectOrientedShowcase::Run(SimpleMemory).0._State_13\.
                            if (\ObjectOrientedShowcase::Run(SimpleMemory).0._State\ = \ObjectOrientedShowcase::Run(SimpleMemory).0._State_16\) then 
                                \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_14\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectOrientedShowcase::Run(SimpleMemory).0._State_17\ => 
                        -- Repeated state of the while loop which was started in state \ObjectOrientedShowcase::Run(SimpleMemory).0._State_14\.
                        -- The while loop's condition:
                        \ObjectOrientedShowcase::Run(SimpleMemory).0.binaryOperationResult.3\ := \ObjectOrientedShowcase::Run(SimpleMemory).0.i\ < to_signed(4, 32);
                        if (\ObjectOrientedShowcase::Run(SimpleMemory).0.binaryOperationResult.3\) then 
                            -- The last invocation for the target state machine finished in the previous state, so need to start the next one in the next state.
                            \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_19\;
                        else 
                            \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_18\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ObjectOrientedShowcase::Run(SimpleMemory).0._State_18\ => 
                        -- State after the while loop which was started in state \ObjectOrientedShowcase::Run(SimpleMemory).0._State_14\.
                        -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.ObjectOrientedShowcase::SumNumberCointainers(Hast.Samples.SampleAssembly.NumberContainer[])
                        \ObjectOrientedShowcase::Run(SimpleMemory).0.ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).numberContainers.parameter.Out.0\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.array\;
                        \ObjectOrientedShowcase::Run(SimpleMemory).0.ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[])._Started.0\ <= true;
                        \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_21\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectOrientedShowcase::Run(SimpleMemory).0._State_19\ => 
                        -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.NumberContainer::IncreaseNumber(System.UInt32)
                        \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32).this.parameter.Out.0\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(\ObjectOrientedShowcase::Run(SimpleMemory).0.i\));
                        \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32).increaseBy.parameter.Out.0\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.array2\(to_integer(to_signed(0, 32))).\Number\;
                        \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32)._Started.0\ <= true;
                        \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_20\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectOrientedShowcase::Run(SimpleMemory).0._State_20\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.NumberContainer::IncreaseNumber(System.UInt32)
                        if (\ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32)._Started.0\ = \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32)._Finished.0\) then 
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32)._Started.0\ <= false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.return.4\ := \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32).return.0\;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.array\(to_integer(\ObjectOrientedShowcase::Run(SimpleMemory).0.i\)) := \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32).this.parameter.In.0\;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.binaryOperationResult.4\ := \ObjectOrientedShowcase::Run(SimpleMemory).0.i\ + to_signed(1, 32);
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.i\ := \ObjectOrientedShowcase::Run(SimpleMemory).0.binaryOperationResult.4\;
                            -- Returning to the repeated state of the while loop which was started in state \ObjectOrientedShowcase::Run(SimpleMemory).0._State_14\ if the loop wasn't exited with a state change.
                            if (\ObjectOrientedShowcase::Run(SimpleMemory).0._State\ = \ObjectOrientedShowcase::Run(SimpleMemory).0._State_20\) then 
                                \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_17\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ObjectOrientedShowcase::Run(SimpleMemory).0._State_21\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.ObjectOrientedShowcase::SumNumberCointainers(Hast.Samples.SampleAssembly.NumberContainer[])
                        if (\ObjectOrientedShowcase::Run(SimpleMemory).0.ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[])._Started.0\ = \ObjectOrientedShowcase::Run(SimpleMemory).0.ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[])._Finished.0\) then 
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[])._Started.0\ <= false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.return.5\ := \ObjectOrientedShowcase::Run(SimpleMemory).0.ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).return.0\;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.array\ := \ObjectOrientedShowcase::Run(SimpleMemory).0.ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).numberContainers.parameter.In.0\;
                            -- Begin SimpleMemory write.
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(to_signed(0, 32), 32);
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.SimpleMemory.WriteEnable\ <= true;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.SimpleMemory.DataOut\ <= ConvertUInt32ToStdLogicVector(\ObjectOrientedShowcase::Run(SimpleMemory).0.return.5\);
                            \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_22\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectOrientedShowcase::Run(SimpleMemory).0._State_22\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \ObjectOrientedShowcase::Run(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                            \ObjectOrientedShowcase::Run(SimpleMemory).0._State\ := \ObjectOrientedShowcase::Run(SimpleMemory).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.Samples.SampleAssembly.ObjectOrientedShowcase::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine end


    -- System.UInt32 Hast.Samples.SampleAssembly.ObjectOrientedShowcase::SumNumberCointainers(Hast.Samples.SampleAssembly.NumberContainer[]).0 state machine start
    \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._StateMachine\: process (\Clock\) 
        Variable \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State\: \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._States\ := \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State_0\;
        Variable \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.numberContainers\: \Hast.Samples.SampleAssembly.NumberContainer_Array\(0 to 3);
        Variable \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.i\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.binaryOperationResult.0\: boolean := false;
        Variable \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.binaryOperationResult.1\: boolean := false;
        Variable \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.binaryOperationResult.2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.binaryOperationResult.3\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._Finished\ <= false;
                \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.return\ <= to_unsigned(0, 32);
                \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State\ := \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State_0\;
                \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.num\ := to_unsigned(0, 32);
                \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.i\ := to_signed(0, 32);
                \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.binaryOperationResult.0\ := false;
                \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.binaryOperationResult.1\ := false;
                \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.binaryOperationResult.2\ := to_unsigned(0, 32);
                \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.binaryOperationResult.3\ := to_signed(0, 32);
            else 
                case \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State\ is 
                    when \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._Started\ = true) then 
                            \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State\ := \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._Started\ = true) then 
                            \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._Finished\ <= true;
                        else 
                            \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._Finished\ <= false;
                            \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State\ := \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.numberContainers.parameter.Out\ <= \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.numberContainers\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State_2\ => 
                        \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.numberContainers\ := \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.numberContainers.parameter.In\;
                        \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.num\ := to_unsigned(0, 32);
                        \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.i\ := to_signed(0, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.binaryOperationResult.0\ := \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.i\ < to_signed(4, 32);
                        if (\ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.binaryOperationResult.0\) then 
                            \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State\ := \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State_3\;
                        else 
                            \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State\ := \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State_3\ => 
                        -- Repeated state of the while loop which was started in state \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State_2\.
                        -- The while loop's condition:
                        \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.binaryOperationResult.1\ := \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.i\ < to_signed(4, 32);
                        if (\ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.binaryOperationResult.1\) then 
                            \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.binaryOperationResult.2\ := \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.num\ + \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.numberContainers\(to_integer(\ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.i\)).\Number\;
                            \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.num\ := \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.binaryOperationResult.2\;
                            \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.binaryOperationResult.3\ := \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.i\ + to_signed(1, 32);
                            \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.i\ := \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.binaryOperationResult.3\;
                        else 
                            \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State\ := \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State_4\ => 
                        -- State after the while loop which was started in state \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State_2\.
                        \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.return\ <= \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.num\;
                        \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State\ := \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.UInt32 Hast.Samples.SampleAssembly.ObjectOrientedShowcase::SumNumberCointainers(Hast.Samples.SampleAssembly.NumberContainer[]).0 state machine end


    -- System.Void Hast.Samples.SampleAssembly.NumberContainer::.ctor().0 state machine start
    \NumberContainer::.ctor().0._StateMachine\: process (\Clock\) 
        Variable \NumberContainer::.ctor().0._State\: \NumberContainer::.ctor().0._States\ := \NumberContainer::.ctor().0._State_0\;
        Variable \NumberContainer::.ctor().0.this\: \Hast.Samples.SampleAssembly.NumberContainer\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \NumberContainer::.ctor().0._Finished\ <= false;
                \NumberContainer::.ctor().0._State\ := \NumberContainer::.ctor().0._State_0\;
            else 
                case \NumberContainer::.ctor().0._State\ is 
                    when \NumberContainer::.ctor().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\NumberContainer::.ctor().0._Started\ = true) then 
                            \NumberContainer::.ctor().0._State\ := \NumberContainer::.ctor().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \NumberContainer::.ctor().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\NumberContainer::.ctor().0._Started\ = true) then 
                            \NumberContainer::.ctor().0._Finished\ <= true;
                        else 
                            \NumberContainer::.ctor().0._Finished\ <= false;
                            \NumberContainer::.ctor().0._State\ := \NumberContainer::.ctor().0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \NumberContainer::.ctor().0.this.parameter.Out\ <= \NumberContainer::.ctor().0.this\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \NumberContainer::.ctor().0._State_2\ => 
                        \NumberContainer::.ctor().0.this\ := \NumberContainer::.ctor().0.this.parameter.In\;
                        \NumberContainer::.ctor().0.this\.\Number\ := to_unsigned(99, 32);
                        \NumberContainer::.ctor().0._State\ := \NumberContainer::.ctor().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.Samples.SampleAssembly.NumberContainer::.ctor().0 state machine end


    -- System.Void Hast.Samples.SampleAssembly.NumberContainer::.ctor(System.UInt32).0 state machine start
    \NumberContainer::.ctor(UInt32).0._StateMachine\: process (\Clock\) 
        Variable \NumberContainer::.ctor(UInt32).0._State\: \NumberContainer::.ctor(UInt32).0._States\ := \NumberContainer::.ctor(UInt32).0._State_0\;
        Variable \NumberContainer::.ctor(UInt32).0.this\: \Hast.Samples.SampleAssembly.NumberContainer\;
        Variable \NumberContainer::.ctor(UInt32).0.number\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \NumberContainer::.ctor(UInt32).0._Finished\ <= false;
                \NumberContainer::.ctor(UInt32).0._State\ := \NumberContainer::.ctor(UInt32).0._State_0\;
                \NumberContainer::.ctor(UInt32).0.number\ := to_unsigned(0, 32);
            else 
                case \NumberContainer::.ctor(UInt32).0._State\ is 
                    when \NumberContainer::.ctor(UInt32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\NumberContainer::.ctor(UInt32).0._Started\ = true) then 
                            \NumberContainer::.ctor(UInt32).0._State\ := \NumberContainer::.ctor(UInt32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \NumberContainer::.ctor(UInt32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\NumberContainer::.ctor(UInt32).0._Started\ = true) then 
                            \NumberContainer::.ctor(UInt32).0._Finished\ <= true;
                        else 
                            \NumberContainer::.ctor(UInt32).0._Finished\ <= false;
                            \NumberContainer::.ctor(UInt32).0._State\ := \NumberContainer::.ctor(UInt32).0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \NumberContainer::.ctor(UInt32).0.this.parameter.Out\ <= \NumberContainer::.ctor(UInt32).0.this\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \NumberContainer::.ctor(UInt32).0._State_2\ => 
                        \NumberContainer::.ctor(UInt32).0.this\ := \NumberContainer::.ctor(UInt32).0.this.parameter.In\;
                        \NumberContainer::.ctor(UInt32).0.number\ := \NumberContainer::.ctor(UInt32).0.number.parameter.In\;
                        \NumberContainer::.ctor(UInt32).0.this\.\Number\ := to_unsigned(99, 32);
                        \NumberContainer::.ctor(UInt32).0.this\.\Number\ := to_unsigned(9, 32);
                        \NumberContainer::.ctor(UInt32).0._State\ := \NumberContainer::.ctor(UInt32).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.Samples.SampleAssembly.NumberContainer::.ctor(System.UInt32).0 state machine end


    -- System.UInt32 Hast.Samples.SampleAssembly.NumberContainer::IncreaseNumber(System.UInt32).0 state machine start
    \NumberContainer::IncreaseNumber(UInt32).0._StateMachine\: process (\Clock\) 
        Variable \NumberContainer::IncreaseNumber(UInt32).0._State\: \NumberContainer::IncreaseNumber(UInt32).0._States\ := \NumberContainer::IncreaseNumber(UInt32).0._State_0\;
        Variable \NumberContainer::IncreaseNumber(UInt32).0.this\: \Hast.Samples.SampleAssembly.NumberContainer\;
        Variable \NumberContainer::IncreaseNumber(UInt32).0.increaseBy\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \NumberContainer::IncreaseNumber(UInt32).0.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \NumberContainer::IncreaseNumber(UInt32).0._Finished\ <= false;
                \NumberContainer::IncreaseNumber(UInt32).0.return\ <= to_unsigned(0, 32);
                \NumberContainer::IncreaseNumber(UInt32).0._State\ := \NumberContainer::IncreaseNumber(UInt32).0._State_0\;
                \NumberContainer::IncreaseNumber(UInt32).0.increaseBy\ := to_unsigned(0, 32);
                \NumberContainer::IncreaseNumber(UInt32).0.binaryOperationResult.0\ := to_unsigned(0, 32);
            else 
                case \NumberContainer::IncreaseNumber(UInt32).0._State\ is 
                    when \NumberContainer::IncreaseNumber(UInt32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\NumberContainer::IncreaseNumber(UInt32).0._Started\ = true) then 
                            \NumberContainer::IncreaseNumber(UInt32).0._State\ := \NumberContainer::IncreaseNumber(UInt32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \NumberContainer::IncreaseNumber(UInt32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\NumberContainer::IncreaseNumber(UInt32).0._Started\ = true) then 
                            \NumberContainer::IncreaseNumber(UInt32).0._Finished\ <= true;
                        else 
                            \NumberContainer::IncreaseNumber(UInt32).0._Finished\ <= false;
                            \NumberContainer::IncreaseNumber(UInt32).0._State\ := \NumberContainer::IncreaseNumber(UInt32).0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \NumberContainer::IncreaseNumber(UInt32).0.this.parameter.Out\ <= \NumberContainer::IncreaseNumber(UInt32).0.this\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \NumberContainer::IncreaseNumber(UInt32).0._State_2\ => 
                        \NumberContainer::IncreaseNumber(UInt32).0.this\ := \NumberContainer::IncreaseNumber(UInt32).0.this.parameter.In\;
                        \NumberContainer::IncreaseNumber(UInt32).0.increaseBy\ := \NumberContainer::IncreaseNumber(UInt32).0.increaseBy.parameter.In\;
                        \NumberContainer::IncreaseNumber(UInt32).0.this\.\WasIncreased\ := True;
                        \NumberContainer::IncreaseNumber(UInt32).0.binaryOperationResult.0\ := \NumberContainer::IncreaseNumber(UInt32).0.this\.\Number\ + \NumberContainer::IncreaseNumber(UInt32).0.increaseBy\;
                        \NumberContainer::IncreaseNumber(UInt32).0.this\.\Number\ := \NumberContainer::IncreaseNumber(UInt32).0.binaryOperationResult.0\;
                        \NumberContainer::IncreaseNumber(UInt32).0.return\ <= \NumberContainer::IncreaseNumber(UInt32).0.this\.\Number\;
                        \NumberContainer::IncreaseNumber(UInt32).0._State\ := \NumberContainer::IncreaseNumber(UInt32).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.UInt32 Hast.Samples.SampleAssembly.NumberContainer::IncreaseNumber(System.UInt32).0 state machine end


    -- System.UInt32 Hast.Samples.SampleAssembly.NumberContainer::get_NumberPlusFive().0 state machine start
    \NumberContainer::get_NumberPlusFive().0._StateMachine\: process (\Clock\) 
        Variable \NumberContainer::get_NumberPlusFive().0._State\: \NumberContainer::get_NumberPlusFive().0._States\ := \NumberContainer::get_NumberPlusFive().0._State_0\;
        Variable \NumberContainer::get_NumberPlusFive().0.this\: \Hast.Samples.SampleAssembly.NumberContainer\;
        Variable \NumberContainer::get_NumberPlusFive().0.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \NumberContainer::get_NumberPlusFive().0._Finished\ <= false;
                \NumberContainer::get_NumberPlusFive().0.return\ <= to_unsigned(0, 32);
                \NumberContainer::get_NumberPlusFive().0._State\ := \NumberContainer::get_NumberPlusFive().0._State_0\;
                \NumberContainer::get_NumberPlusFive().0.binaryOperationResult.0\ := to_unsigned(0, 32);
            else 
                case \NumberContainer::get_NumberPlusFive().0._State\ is 
                    when \NumberContainer::get_NumberPlusFive().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\NumberContainer::get_NumberPlusFive().0._Started\ = true) then 
                            \NumberContainer::get_NumberPlusFive().0._State\ := \NumberContainer::get_NumberPlusFive().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \NumberContainer::get_NumberPlusFive().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\NumberContainer::get_NumberPlusFive().0._Started\ = true) then 
                            \NumberContainer::get_NumberPlusFive().0._Finished\ <= true;
                        else 
                            \NumberContainer::get_NumberPlusFive().0._Finished\ <= false;
                            \NumberContainer::get_NumberPlusFive().0._State\ := \NumberContainer::get_NumberPlusFive().0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \NumberContainer::get_NumberPlusFive().0.this.parameter.Out\ <= \NumberContainer::get_NumberPlusFive().0.this\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \NumberContainer::get_NumberPlusFive().0._State_2\ => 
                        \NumberContainer::get_NumberPlusFive().0.this\ := \NumberContainer::get_NumberPlusFive().0.this.parameter.In\;
                        \NumberContainer::get_NumberPlusFive().0.binaryOperationResult.0\ := \NumberContainer::get_NumberPlusFive().0.this\.\Number\ + to_unsigned(5, 32);
                        \NumberContainer::get_NumberPlusFive().0.return\ <= \NumberContainer::get_NumberPlusFive().0.binaryOperationResult.0\;
                        \NumberContainer::get_NumberPlusFive().0._State\ := \NumberContainer::get_NumberPlusFive().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.UInt32 Hast.Samples.SampleAssembly.NumberContainer::get_NumberPlusFive().0 state machine end


    -- System.Void Hast.Samples.SampleAssembly.NumberContainer::set_NumberPlusFive(System.UInt32).0 state machine start
    \NumberContainer::set_NumberPlusFive(UInt32).0._StateMachine\: process (\Clock\) 
        Variable \NumberContainer::set_NumberPlusFive(UInt32).0._State\: \NumberContainer::set_NumberPlusFive(UInt32).0._States\ := \NumberContainer::set_NumberPlusFive(UInt32).0._State_0\;
        Variable \NumberContainer::set_NumberPlusFive(UInt32).0.this\: \Hast.Samples.SampleAssembly.NumberContainer\;
        Variable \NumberContainer::set_NumberPlusFive(UInt32).0.value\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \NumberContainer::set_NumberPlusFive(UInt32).0.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \NumberContainer::set_NumberPlusFive(UInt32).0._Finished\ <= false;
                \NumberContainer::set_NumberPlusFive(UInt32).0._State\ := \NumberContainer::set_NumberPlusFive(UInt32).0._State_0\;
                \NumberContainer::set_NumberPlusFive(UInt32).0.value\ := to_unsigned(0, 32);
                \NumberContainer::set_NumberPlusFive(UInt32).0.binaryOperationResult.0\ := to_unsigned(0, 32);
            else 
                case \NumberContainer::set_NumberPlusFive(UInt32).0._State\ is 
                    when \NumberContainer::set_NumberPlusFive(UInt32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\NumberContainer::set_NumberPlusFive(UInt32).0._Started\ = true) then 
                            \NumberContainer::set_NumberPlusFive(UInt32).0._State\ := \NumberContainer::set_NumberPlusFive(UInt32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \NumberContainer::set_NumberPlusFive(UInt32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\NumberContainer::set_NumberPlusFive(UInt32).0._Started\ = true) then 
                            \NumberContainer::set_NumberPlusFive(UInt32).0._Finished\ <= true;
                        else 
                            \NumberContainer::set_NumberPlusFive(UInt32).0._Finished\ <= false;
                            \NumberContainer::set_NumberPlusFive(UInt32).0._State\ := \NumberContainer::set_NumberPlusFive(UInt32).0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \NumberContainer::set_NumberPlusFive(UInt32).0.this.parameter.Out\ <= \NumberContainer::set_NumberPlusFive(UInt32).0.this\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \NumberContainer::set_NumberPlusFive(UInt32).0._State_2\ => 
                        \NumberContainer::set_NumberPlusFive(UInt32).0.this\ := \NumberContainer::set_NumberPlusFive(UInt32).0.this.parameter.In\;
                        \NumberContainer::set_NumberPlusFive(UInt32).0.value\ := \NumberContainer::set_NumberPlusFive(UInt32).0.value.parameter.In\;
                        \NumberContainer::set_NumberPlusFive(UInt32).0.binaryOperationResult.0\ := \NumberContainer::set_NumberPlusFive(UInt32).0.value\ - to_unsigned(5, 32);
                        \NumberContainer::set_NumberPlusFive(UInt32).0.this\.\Number\ := \NumberContainer::set_NumberPlusFive(UInt32).0.binaryOperationResult.0\;
                        \NumberContainer::set_NumberPlusFive(UInt32).0._State\ := \NumberContainer::set_NumberPlusFive(UInt32).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.Samples.SampleAssembly.NumberContainer::set_NumberPlusFive(System.UInt32).0 state machine end


    -- System.Void Hast.Samples.SampleAssembly.MemoryContainer::.ctor(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine start
    \MemoryContainer::.ctor(SimpleMemory).0._StateMachine\: process (\Clock\) 
        Variable \MemoryContainer::.ctor(SimpleMemory).0._State\: \MemoryContainer::.ctor(SimpleMemory).0._States\ := \MemoryContainer::.ctor(SimpleMemory).0._State_0\;
        Variable \MemoryContainer::.ctor(SimpleMemory).0.this\: \Hast.Samples.SampleAssembly.MemoryContainer\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \MemoryContainer::.ctor(SimpleMemory).0._Finished\ <= false;
                \MemoryContainer::.ctor(SimpleMemory).0._State\ := \MemoryContainer::.ctor(SimpleMemory).0._State_0\;
            else 
                case \MemoryContainer::.ctor(SimpleMemory).0._State\ is 
                    when \MemoryContainer::.ctor(SimpleMemory).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\MemoryContainer::.ctor(SimpleMemory).0._Started\ = true) then 
                            \MemoryContainer::.ctor(SimpleMemory).0._State\ := \MemoryContainer::.ctor(SimpleMemory).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \MemoryContainer::.ctor(SimpleMemory).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\MemoryContainer::.ctor(SimpleMemory).0._Started\ = true) then 
                            \MemoryContainer::.ctor(SimpleMemory).0._Finished\ <= true;
                        else 
                            \MemoryContainer::.ctor(SimpleMemory).0._Finished\ <= false;
                            \MemoryContainer::.ctor(SimpleMemory).0._State\ := \MemoryContainer::.ctor(SimpleMemory).0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \MemoryContainer::.ctor(SimpleMemory).0.this.parameter.Out\ <= \MemoryContainer::.ctor(SimpleMemory).0.this\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \MemoryContainer::.ctor(SimpleMemory).0._State_2\ => 
                        \MemoryContainer::.ctor(SimpleMemory).0.this\ := \MemoryContainer::.ctor(SimpleMemory).0.this.parameter.In\;
                        \MemoryContainer::.ctor(SimpleMemory).0._State\ := \MemoryContainer::.ctor(SimpleMemory).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.Samples.SampleAssembly.MemoryContainer::.ctor(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine end


    -- System.UInt32 Hast.Samples.SampleAssembly.MemoryContainer::GetInput().0 state machine start
    \MemoryContainer::GetInput().0._StateMachine\: process (\Clock\) 
        Variable \MemoryContainer::GetInput().0._State\: \MemoryContainer::GetInput().0._States\ := \MemoryContainer::GetInput().0._State_0\;
        Variable \MemoryContainer::GetInput().0.this\: \Hast.Samples.SampleAssembly.MemoryContainer\;
        Variable \MemoryContainer::GetInput().0.dataIn.0\: std_logic_vector(31 downto 0);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \MemoryContainer::GetInput().0._Finished\ <= false;
                \MemoryContainer::GetInput().0.return\ <= to_unsigned(0, 32);
                \MemoryContainer::GetInput().0.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \MemoryContainer::GetInput().0.SimpleMemory.ReadEnable\ <= false;
                \MemoryContainer::GetInput().0.SimpleMemory.WriteEnable\ <= false;
                \MemoryContainer::GetInput().0._State\ := \MemoryContainer::GetInput().0._State_0\;
            else 
                case \MemoryContainer::GetInput().0._State\ is 
                    when \MemoryContainer::GetInput().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\MemoryContainer::GetInput().0._Started\ = true) then 
                            \MemoryContainer::GetInput().0._State\ := \MemoryContainer::GetInput().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \MemoryContainer::GetInput().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\MemoryContainer::GetInput().0._Started\ = true) then 
                            \MemoryContainer::GetInput().0._Finished\ <= true;
                        else 
                            \MemoryContainer::GetInput().0._Finished\ <= false;
                            \MemoryContainer::GetInput().0._State\ := \MemoryContainer::GetInput().0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \MemoryContainer::GetInput().0.this.parameter.Out\ <= \MemoryContainer::GetInput().0.this\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \MemoryContainer::GetInput().0._State_2\ => 
                        \MemoryContainer::GetInput().0.this\ := \MemoryContainer::GetInput().0.this.parameter.In\;
                        -- Begin SimpleMemory read.
                        \MemoryContainer::GetInput().0.SimpleMemory.CellIndex\ <= resize(to_signed(0, 32), 32);
                        \MemoryContainer::GetInput().0.SimpleMemory.ReadEnable\ <= true;
                        \MemoryContainer::GetInput().0._State\ := \MemoryContainer::GetInput().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \MemoryContainer::GetInput().0._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \MemoryContainer::GetInput().0.SimpleMemory.ReadEnable\ <= false;
                            \MemoryContainer::GetInput().0.dataIn.0\ := \DataIn\;
                            \MemoryContainer::GetInput().0.return\ <= ConvertStdLogicVectorToUInt32(\MemoryContainer::GetInput().0.dataIn.0\);
                            \MemoryContainer::GetInput().0._State\ := \MemoryContainer::GetInput().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.UInt32 Hast.Samples.SampleAssembly.MemoryContainer::GetInput().0 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32).0 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.numberObject\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.num2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.num3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.flag\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.result\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.1\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.2\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.4\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.5\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.return\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.numberObject\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.num\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.num2\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.num3\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.flag\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.result\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.0\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.1\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.2\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.3\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.4\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.5\ := to_unsigned(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.numberObject.parameter.In\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.return\ <= True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.num3\;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32).0 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32).1 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.numberObject\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.num2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.num3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.flag\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.result\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.1\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.2\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.4\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.5\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.return\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.numberObject\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.num\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.num2\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.num3\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.flag\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.result\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.0\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.1\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.2\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.3\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.4\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.5\ := to_unsigned(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.numberObject.parameter.In\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.return\ <= True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.num3\;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32).1 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32).2 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.numberObject\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.num2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.num3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.flag\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.result\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.1\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.2\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.4\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.5\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.return\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.numberObject\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.num\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.num2\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.num3\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.flag\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.result\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.0\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.1\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.2\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.3\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.4\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.5\ := to_unsigned(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.numberObject.parameter.In\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.return\ <= True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.num3\;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32).2 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32).3 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.numberObject\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.num2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.num3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.flag\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.result\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.1\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.2\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.4\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.5\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.return\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.numberObject\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.num\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.num2\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.num3\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.flag\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.result\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.0\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.1\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.2\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.3\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.4\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.5\ := to_unsigned(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.numberObject.parameter.In\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.return\ <= True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.num3\;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32).3 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32).4 state machine start
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State\: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._States\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_0\;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.numberObject\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.num2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.num3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.flag\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.result\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.1\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.2\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.4\: boolean := false;
        Variable \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.5\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._Finished\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.return\ <= false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_0\;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.numberObject\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.num\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.num2\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.num3\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.flag\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.result\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.0\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.1\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.2\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.3\ := to_unsigned(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.4\ := false;
                \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.5\ := to_unsigned(0, 32);
            else 
                case \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State\ is 
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._Started\ = true) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._Finished\ <= true;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._Finished\ <= false;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_2\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.numberObject\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.numberObject.parameter.In\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.num\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.numberObject\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.num\ / to_unsigned(2, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.num2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.0\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.num3\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.1\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.1\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_3\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.2\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.num3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.num2\;
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.2\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_5\;
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_2\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.result\ := True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.return\ <= True;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_6\;
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.num\ mod \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.num3\;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_6\ => 
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.4\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.flag\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_8\ and ends in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_7\.

                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.flag\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.5\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.num3\ + to_unsigned(1, 32);
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.num3\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_7\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_6\.
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.result\ := False;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.return\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.result\;
                        \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_6\.
                        if (\PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State\ = \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_8\) then 
                            \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State\ := \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32).4 state machine end


    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumber(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine start
    \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State\: \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._States\ := \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_0\;
        Variable \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.number\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.dataIn.0\: std_logic_vector(31 downto 0);
        Variable \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.return.0\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Finished\ <= false;
                \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).number.parameter.Out.0\ <= to_unsigned(0, 32);
                \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\ <= false;
                \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_0\;
                \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.number\ := to_unsigned(0, 32);
                \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.return.0\ := false;
            else 
                case \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State\ is 
                    when \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Started\ = true) then 
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Started\ = true) then 
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Finished\ <= true;
                        else 
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Finished\ <= false;
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_2\ => 
                        -- Begin SimpleMemory read.
                        \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(to_signed(0, 32), 32);
                        \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.ReadEnable\ <= true;
                        \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.dataIn.0\ := \DataIn\;
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.number\ := ConvertStdLogicVectorToUInt32(\PrimeCalculator::IsPrimeNumber(SimpleMemory).0.dataIn.0\);
                            -- Starting state machine invocation for the following method: System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberInternal(System.UInt32)
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).number.parameter.Out.0\ <= \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.number\;
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\ <= true;
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberInternal(System.UInt32)
                        if (\PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\ = \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\) then 
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\ <= false;
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.return.0\ := \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).return.0\;
                            -- Begin SimpleMemory write.
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(to_signed(0, 32), 32);
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.WriteEnable\ <= true;
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.DataOut\ <= ConvertBooleanToStdLogicVector(\PrimeCalculator::IsPrimeNumber(SimpleMemory).0.return.0\);
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_5\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumber(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine end


    -- System.Threading.Tasks.Task Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberAsync(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine start
    \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State\: \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._States\ := \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_0\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._Finished\ <= false;
                \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\ <= false;
                \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_0\;
            else 
                case \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State\ is 
                    when \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._Started\ = true) then 
                            \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._Started\ = true) then 
                            \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._Finished\ <= true;
                        else 
                            \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._Finished\ <= false;
                            \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_2\ => 
                        -- Starting state machine invocation for the following method: System.Void Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumber(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory)
                        \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\ <= true;
                        \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumber(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory)
                        if (\PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\ = \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\) then 
                            \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\ <= false;
                            \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State\ := \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Threading.Tasks.Task Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberAsync(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine end


    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ArePrimeNumbers(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine start
    \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\: \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._States\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_0\;
        Variable \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.number\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.dataIn.0\: std_logic_vector(31 downto 0);
        Variable \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.0\: boolean := false;
        Variable \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.1\: boolean := false;
        Variable \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.dataIn.1\: std_logic_vector(31 downto 0);
        Variable \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.3\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.return.0\: boolean := false;
        Variable \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.4\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._Finished\ <= false;
                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).number.parameter.Out.0\ <= to_unsigned(0, 32);
                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\ <= false;
                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_0\;
                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num\ := to_unsigned(0, 32);
                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num2\ := to_signed(0, 32);
                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.number\ := to_unsigned(0, 32);
                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.0\ := false;
                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.1\ := false;
                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.2\ := to_signed(0, 32);
                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.3\ := to_signed(0, 32);
                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.return.0\ := false;
                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.4\ := to_signed(0, 32);
            else 
                case \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ is 
                    when \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._Started\ = true) then 
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._Started\ = true) then 
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._Finished\ <= true;
                        else 
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._Finished\ <= false;
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_2\ => 
                        -- Begin SimpleMemory read.
                        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(to_signed(0, 32), 32);
                        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ <= true;
                        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.dataIn.0\ := \DataIn\;
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num\ := ConvertStdLogicVectorToUInt32(\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.dataIn.0\);
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num2\ := to_signed(0, 32);
                            -- Starting a while loop.
                            -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.0\ := resize(\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num2\, 64) < signed((resize(\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num\, 64)));
                            if (\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.0\) then 
                                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_4\;
                            else 
                                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_5\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_4\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_3\.
                        -- The while loop's condition:
                        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.1\ := resize(\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num2\, 64) < signed((resize(\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num\, 64)));
                        if (\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.1\) then 
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.2\ := to_signed(1, 32) + \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num2\;
                            -- Begin SimpleMemory read.
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.2\, 32);
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ <= true;
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_6\;
                        else 
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_5\ => 
                        -- State after the while loop which was started in state \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_3\.
                        \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_6\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.dataIn.1\ := \DataIn\;
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.number\ := ConvertStdLogicVectorToUInt32(\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.dataIn.1\);
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.3\ := to_signed(1, 32) + \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num2\;
                            -- Starting state machine invocation for the following method: System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberInternal(System.UInt32)
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).number.parameter.Out.0\ <= \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.number\;
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\ <= true;
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_7\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberInternal(System.UInt32)
                        if (\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\ = \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\) then 
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\ <= false;
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.return.0\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).return.0\;
                            -- Begin SimpleMemory write.
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.3\, 32);
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ <= true;
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.DataOut\ <= ConvertBooleanToStdLogicVector(\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.return.0\);
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_8\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.4\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num2\ + to_signed(1, 32);
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.num2\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.binaryOperationResult.4\;
                            -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_3\ if the loop wasn't exited with a state change.
                            if (\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ = \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_8\) then 
                                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._State_4\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ArePrimeNumbers(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine end


    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine start
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\: \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._States\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_0\;
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\: \boolean_Array\(0 to 29) := (others => false);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.i\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.arg_5D_1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.j\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.dataIn.0\: std_logic_vector(31 downto 0);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.0\: boolean := false;
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.1\: boolean := false;
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.2\: boolean := false;
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.3\: boolean := false;
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.4\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.5\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.dataIn.1\: std_logic_vector(31 downto 0);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).invocationIndex\: integer range 0 to 4 := 0;
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.6\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.return.0\: boolean := false;
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.return.1\: boolean := false;
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.return.2\: boolean := false;
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.return.3\: boolean := false;
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.return.4\: boolean := false;
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.7\: boolean := false;
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.8\: boolean := false;
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.9\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.10\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.11\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.12\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._Finished\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).numberObject.parameter.Out.0\ <= to_unsigned(0, 32);
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.0\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).numberObject.parameter.Out.1\ <= to_unsigned(0, 32);
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.1\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).numberObject.parameter.Out.2\ <= to_unsigned(0, 32);
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.2\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).numberObject.parameter.Out.3\ <= to_unsigned(0, 32);
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.3\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).numberObject.parameter.Out.4\ <= to_unsigned(0, 32);
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.4\ <= false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_0\;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num\ := to_unsigned(0, 32);
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\ := (others => false);
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num2\ := to_signed(0, 32);
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.i\ := to_signed(0, 32);
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\ := to_unsigned(0, 32);
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.arg_5D_1\ := to_signed(0, 32);
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.j\ := to_signed(0, 32);
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.0\ := false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.1\ := false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.2\ := false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.3\ := false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.4\ := to_signed(0, 32);
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.5\ := to_signed(0, 32);
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).invocationIndex\ := 0;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.6\ := to_signed(0, 32);
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.return.0\ := false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.return.1\ := false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.return.2\ := false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.return.3\ := false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.return.4\ := false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.7\ := false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.8\ := false;
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.9\ := to_signed(0, 32);
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.10\ := to_signed(0, 32);
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.11\ := to_signed(0, 32);
                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.12\ := to_signed(0, 32);
            else 
                case \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ is 
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._Started\ = true) then 
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._Started\ = true) then 
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._Finished\ <= true;
                        else 
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._Finished\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_2\ => 
                        -- Begin SimpleMemory read.
                        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(to_signed(0, 32), 32);
                        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ <= true;
                        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.dataIn.0\ := \DataIn\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num\ := ConvertStdLogicVectorToUInt32(\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.dataIn.0\);
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\ := (others => false);
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num2\ := to_signed(0, 32);
                            -- Starting a while loop.
                            -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.0\ := resize(\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num2\, 64) < signed((resize(\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num\, 64)));
                            if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.0\) then 
                                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_4\;
                            else 
                                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_5\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_4\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_3\.
                        -- The while loop's condition:
                        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.1\ := resize(\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num2\, 64) < signed((resize(\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num\, 64)));
                        if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.1\) then 
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.i\ := to_signed(0, 32);
                            -- Starting a while loop.
                            -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.2\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.i\ < to_signed(30, 32);
                            if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.2\) then 
                                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_6\;
                            else 
                                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_7\;
                            end if;
                        else 
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_5\ => 
                        -- State after the while loop which was started in state \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_3\.
                        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_6\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_4\.
                        -- The while loop's condition:
                        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.3\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.i\ < to_signed(30, 32);
                        if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.3\) then 
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.4\ := to_signed(1, 32) + \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num2\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.5\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.4\ + \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.i\;
                            -- Begin SimpleMemory read.
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.5\, 32);
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ <= true;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_8\;
                        else 
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_7\ => 
                        -- State after the while loop which was started in state \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_4\.
                        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_9\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_8\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.dataIn.1\ := \DataIn\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\ := ConvertStdLogicVectorToUInt32(\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.dataIn.1\);
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.arg_5D_1\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.i\;
                            -- Starting state machine invocation for the following method: System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32)
                            case \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).invocationIndex\ is 
                                when 0 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).numberObject.parameter.Out.0\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.0\ <= true;
                                when 1 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).numberObject.parameter.Out.1\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.1\ <= true;
                                when 2 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).numberObject.parameter.Out.2\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.2\ <= true;
                                when 3 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).numberObject.parameter.Out.3\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.3\ <= true;
                                when 4 => 
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).numberObject.parameter.Out.4\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num3\;
                                    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.4\ <= true;
                            end case;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).invocationIndex\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).invocationIndex\ + 1;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.6\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.i\ + to_signed(1, 32);
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.i\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.6\;
                            -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_4\ if the loop wasn't exited with a state change.
                            if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_8\) then 
                                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_6\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_9\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32)
                        if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.1\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Finished.1\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.2\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Finished.2\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.3\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Finished.3\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.4\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Finished.4\ and \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.0\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Finished.0\) then 
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.0\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.1\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.2\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.3\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.4\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).invocationIndex\ := 0;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.return.0\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).return.0\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.return.1\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).return.1\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.return.2\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).return.2\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.return.3\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).return.3\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.return.4\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).return.4\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(0) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.return.0\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(1) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.return.1\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(2) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.return.2\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(3) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.return.3\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(4) := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.return.4\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.j\ := to_signed(0, 32);
                            -- Starting a while loop.
                            -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.7\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.j\ < to_signed(30, 32);
                            if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.7\) then 
                                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_10\;
                            else 
                                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_11\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_10\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_9\.
                        -- The while loop's condition:
                        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.8\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.j\ < to_signed(30, 32);
                        if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.8\) then 
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.9\ := to_signed(1, 32) + \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num2\;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.10\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.9\ + \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.j\;
                            -- Begin SimpleMemory write.
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.10\, 32);
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ <= true;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.DataOut\ <= ConvertBooleanToStdLogicVector(\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.array\(to_integer(\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.j\)));
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_12\;
                        else 
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_11\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_11\ => 
                        -- State after the while loop which was started in state \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_9\.
                        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.12\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num2\ + to_signed(30, 32);
                        \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.num2\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.12\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_3\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_11\) then 
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_12\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.11\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.j\ + to_signed(1, 32);
                            \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.j\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.binaryOperationResult.11\;
                            -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_9\ if the loop wasn't exited with a state change.
                            if (\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ = \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_12\) then 
                                \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State\ := \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._State_10\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine end


    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberInternal(System.UInt32).0 state machine start
    \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._StateMachine\: process (\Clock\) 
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\: \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._States\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_0\;
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.number\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.flag\: boolean := false;
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.result\: boolean := false;
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.1\: boolean := false;
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.2\: boolean := false;
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.4\: boolean := false;
        Variable \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.5\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Finished\ <= false;
                \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.return\ <= false;
                \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_0\;
                \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.number\ := to_unsigned(0, 32);
                \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num\ := to_unsigned(0, 32);
                \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num2\ := to_unsigned(0, 32);
                \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.flag\ := false;
                \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.result\ := false;
                \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.0\ := to_unsigned(0, 32);
                \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.1\ := false;
                \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.2\ := false;
                \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.3\ := to_unsigned(0, 32);
                \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.4\ := false;
                \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.5\ := to_unsigned(0, 32);
            else 
                case \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ is 
                    when \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Started\ = true) then 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Started\ = true) then 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Finished\ <= true;
                        else 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Finished\ <= false;
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_2\ => 
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.number\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.number.parameter.In\;
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.0\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.number\ / to_unsigned(2, 32);
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.0\;
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num2\ := to_unsigned(2, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.1\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num2\ <= \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num\;
                        if (\PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.1\) then 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_3\;
                        else 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_3\ => 
                        -- Repeated state of the while loop which was started in state \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_2\.
                        -- The while loop's condition:
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.2\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num2\ <= \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num\;
                        if (\PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.2\) then 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_5\;
                        else 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_4\ => 
                        -- State after the while loop which was started in state \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_2\.
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.result\ := True;
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.return\ <= True;
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_5\ => 
                        -- Waiting for the result to appear in \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.3\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\PrimeCalculator::IsPrimeNumberInternal(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_6\;
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.3\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.number\ mod \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num2\;
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_6\ => 
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.4\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.3\ = to_unsigned(0, 32);
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.flag\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.4\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_8\ and ends in state \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_8\.
                        --     * Execution after either branch will continue in the following state: \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_7\.

                        if (\PrimeCalculator::IsPrimeNumberInternal(UInt32).0.flag\) then 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_8\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_7\ => 
                        -- State after the if-else which was started in state \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_6\.
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.5\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num2\ + to_unsigned(1, 32);
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.num2\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_2\ if the loop wasn't exited with a state change.
                        if (\PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ = \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_7\) then 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_8\ => 
                        -- True branch of the if-else started in state \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_6\.
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.result\ := False;
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.return\ <= \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.result\;
                        \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_1\;
                        -- Going to the state after the if-else which was started in state \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_6\.
                        if (\PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ = \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_8\) then 
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State\ := \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberInternal(System.UInt32).0 state machine end


    -- System.Void Hast.Samples.SampleAssembly.RecursiveAlgorithms::CalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine start
    \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._StateMachine\: process (\Clock\) 
        Variable \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State\: \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._States\ := \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State_0\;
        Variable \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.number\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.dataIn.0\: std_logic_vector(31 downto 0);
        Variable \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._Finished\ <= false;
                \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\ <= to_signed(0, 16);
                \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= false;
                \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State\ := \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State_0\;
                \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.number\ := to_signed(0, 16);
                \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.return.0\ := to_unsigned(0, 32);
            else 
                case \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State\ is 
                    when \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._Started\ = true) then 
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State\ := \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._Started\ = true) then 
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._Finished\ <= true;
                        else 
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._Finished\ <= false;
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State\ := \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State_2\ => 
                        -- Begin SimpleMemory write.
                        \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                        \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.WriteEnable\ <= true;
                        \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.DataOut\ <= ConvertUInt32ToStdLogicVector(to_unsigned(1, 32));
                        \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State\ := \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                            -- Begin SimpleMemory read.
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(to_signed(0, 32), 32);
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.ReadEnable\ <= true;
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State\ := \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State_4\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.dataIn.0\ := \DataIn\;
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.number\ := resize(ConvertStdLogicVectorToInt32(\RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.dataIn.0\), 16);
                            -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\ <= \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.number\;
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= true;
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State\ := \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        if (\RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ = \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\) then 
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= false;
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.return.0\ := \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\;
                            -- Begin SimpleMemory write.
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(to_signed(0, 32), 32);
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.WriteEnable\ <= true;
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.DataOut\ <= ConvertUInt32ToStdLogicVector(\RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.return.0\);
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State\ := \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State_6\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State\ := \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.Samples.SampleAssembly.RecursiveAlgorithms::CalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine end


    -- System.Void Hast.Samples.SampleAssembly.RecursiveAlgorithms::CalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine start
    \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._StateMachine\: process (\Clock\) 
        Variable \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State\: \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._States\ := \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State_0\;
        Variable \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.number\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.dataIn.0\: std_logic_vector(31 downto 0);
        Variable \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._Finished\ <= false;
                \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\ <= to_signed(0, 16);
                \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ <= false;
                \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State\ := \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State_0\;
                \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.number\ := to_signed(0, 16);
                \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.return.0\ := to_unsigned(0, 32);
            else 
                case \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State\ is 
                    when \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._Started\ = true) then 
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State\ := \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._Started\ = true) then 
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._Finished\ <= true;
                        else 
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._Finished\ <= false;
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State\ := \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State_2\ => 
                        -- Begin SimpleMemory write.
                        \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                        \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.WriteEnable\ <= true;
                        \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.DataOut\ <= ConvertUInt32ToStdLogicVector(to_unsigned(1, 32));
                        \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State\ := \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                            -- Begin SimpleMemory read.
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(to_signed(0, 32), 32);
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.ReadEnable\ <= true;
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State\ := \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State_4\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.dataIn.0\ := \DataIn\;
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.number\ := resize(ConvertStdLogicVectorToInt32(\RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.dataIn.0\), 16);
                            -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\ <= \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.number\;
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ <= true;
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State\ := \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        if (\RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ = \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\) then 
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ <= false;
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.return.0\ := \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\;
                            -- Begin SimpleMemory write.
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(to_signed(0, 32), 32);
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.WriteEnable\ <= true;
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.DataOut\ <= ConvertUInt32ToStdLogicVector(\RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.return.0\);
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State\ := \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State_6\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State\ := \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.Samples.SampleAssembly.RecursiveAlgorithms::CalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).0 state machine start
    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._StateMachine\: process (\Clock\) 
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State\: \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._States\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_0\;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.number\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.flag\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.result\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.dataIn.0\: std_logic_vector(31 downto 0);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.1\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.2\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.3\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.4\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.5\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.return.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.6\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Finished\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.return\ <= to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.SimpleMemory.ReadEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.SimpleMemory.WriteEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\ <= to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_0\;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.number\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.flag\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.result\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.1\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.2\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.3\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.4\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.return.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.5\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.return.1\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.6\ := to_unsigned(0, 32);
            else 
                case \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State\ is 
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Finished\ <= true;
                        else 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Finished\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_2\ => 
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.number\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.number.parameter.In\;
                        -- Begin SimpleMemory read.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.SimpleMemory.ReadEnable\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.SimpleMemory.ReadEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.dataIn.0\ := \DataIn\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.0\ := ConvertStdLogicVectorToUInt32(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.dataIn.0\) + to_unsigned(1, 32);
                            -- Begin SimpleMemory write.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.SimpleMemory.WriteEnable\ <= true;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.SimpleMemory.DataOut\ <= ConvertUInt32ToStdLogicVector(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.0\);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_4\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.SimpleMemory.WriteEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.1\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.number\ = to_signed(0, 16);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.2\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.number\ = to_signed(1, 16);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.3\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.1\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.2\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.flag\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.3\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_6\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_6\.
                            --     * The false branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_7\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_11\.
                            --     * Execution after either branch will continue in the following state: \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_5\.

                            if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.flag\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_6\;
                            else 
                                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_7\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_5\ => 
                        -- State after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.return\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.result\;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_6\ => 
                        -- True branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.result\ := resize(unsigned(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.number\), 32);
                        -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_4\.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_6\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_7\ => 
                        -- False branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.4\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.number\ - to_signed(2, 16);
                        -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.4\;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_8\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_8\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.return.0\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.5\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.number\ - to_signed(1, 16);
                            -- The last invocation for the target state machine just finished, so need to start the next one in a later state.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_9\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_9\ => 
                        -- This state was just added to leave time for the invocation proxy to register that the previous invocation finished.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_10\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_10\ => 
                        -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.5\;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_11\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_11\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.return.1\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.6\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.return.0\ + \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.return.1\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.result\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.binaryOperationResult.6\;
                            -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_4\.
                            if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_11\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._State_5\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).0 state machine end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).1 state machine start
    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._StateMachine\: process (\Clock\) 
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State\: \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._States\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_0\;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.number\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.flag\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.result\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.dataIn.0\: std_logic_vector(31 downto 0);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.1\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.2\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.3\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.4\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.5\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.return.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.6\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Finished\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.return\ <= to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.SimpleMemory.ReadEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.SimpleMemory.WriteEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\ <= to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_0\;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.number\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.flag\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.result\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.1\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.2\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.3\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.4\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.return.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.5\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.return.1\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.6\ := to_unsigned(0, 32);
            else 
                case \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State\ is 
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Finished\ <= true;
                        else 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Finished\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_2\ => 
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.number\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.number.parameter.In\;
                        -- Begin SimpleMemory read.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.SimpleMemory.ReadEnable\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.SimpleMemory.ReadEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.dataIn.0\ := \DataIn\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.0\ := ConvertStdLogicVectorToUInt32(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.dataIn.0\) + to_unsigned(1, 32);
                            -- Begin SimpleMemory write.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.SimpleMemory.WriteEnable\ <= true;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.SimpleMemory.DataOut\ <= ConvertUInt32ToStdLogicVector(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.0\);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_4\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.SimpleMemory.WriteEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.1\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.number\ = to_signed(0, 16);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.2\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.number\ = to_signed(1, 16);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.3\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.1\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.2\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.flag\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.3\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_6\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_6\.
                            --     * The false branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_7\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_11\.
                            --     * Execution after either branch will continue in the following state: \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_5\.

                            if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.flag\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_6\;
                            else 
                                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_7\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_5\ => 
                        -- State after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.return\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.result\;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_6\ => 
                        -- True branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.result\ := resize(unsigned(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.number\), 32);
                        -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_4\.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_6\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_7\ => 
                        -- False branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.4\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.number\ - to_signed(2, 16);
                        -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.4\;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_8\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_8\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.return.0\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.5\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.number\ - to_signed(1, 16);
                            -- The last invocation for the target state machine just finished, so need to start the next one in a later state.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_9\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_9\ => 
                        -- This state was just added to leave time for the invocation proxy to register that the previous invocation finished.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_10\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_10\ => 
                        -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.5\;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_11\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_11\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.return.1\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.6\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.return.0\ + \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.return.1\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.result\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.binaryOperationResult.6\;
                            -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_4\.
                            if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_11\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._State_5\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).1 state machine end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).2 state machine start
    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._StateMachine\: process (\Clock\) 
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State\: \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._States\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_0\;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.number\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.flag\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.result\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.dataIn.0\: std_logic_vector(31 downto 0);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.1\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.2\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.3\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.4\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.5\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.return.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.6\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Finished\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.return\ <= to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.SimpleMemory.ReadEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.SimpleMemory.WriteEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\ <= to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_0\;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.number\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.flag\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.result\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.1\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.2\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.3\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.4\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.return.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.5\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.return.1\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.6\ := to_unsigned(0, 32);
            else 
                case \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State\ is 
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Finished\ <= true;
                        else 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Finished\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_2\ => 
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.number\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.number.parameter.In\;
                        -- Begin SimpleMemory read.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.SimpleMemory.ReadEnable\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.SimpleMemory.ReadEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.dataIn.0\ := \DataIn\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.0\ := ConvertStdLogicVectorToUInt32(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.dataIn.0\) + to_unsigned(1, 32);
                            -- Begin SimpleMemory write.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.SimpleMemory.WriteEnable\ <= true;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.SimpleMemory.DataOut\ <= ConvertUInt32ToStdLogicVector(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.0\);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_4\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.SimpleMemory.WriteEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.1\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.number\ = to_signed(0, 16);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.2\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.number\ = to_signed(1, 16);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.3\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.1\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.2\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.flag\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.3\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_6\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_6\.
                            --     * The false branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_7\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_11\.
                            --     * Execution after either branch will continue in the following state: \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_5\.

                            if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.flag\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_6\;
                            else 
                                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_7\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_5\ => 
                        -- State after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.return\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.result\;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_6\ => 
                        -- True branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.result\ := resize(unsigned(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.number\), 32);
                        -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_4\.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_6\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_7\ => 
                        -- False branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.4\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.number\ - to_signed(2, 16);
                        -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.4\;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_8\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_8\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.return.0\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.5\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.number\ - to_signed(1, 16);
                            -- The last invocation for the target state machine just finished, so need to start the next one in a later state.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_9\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_9\ => 
                        -- This state was just added to leave time for the invocation proxy to register that the previous invocation finished.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_10\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_10\ => 
                        -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.5\;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_11\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_11\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.return.1\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.6\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.return.0\ + \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.return.1\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.result\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.binaryOperationResult.6\;
                            -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_4\.
                            if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_11\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._State_5\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).2 state machine end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).3 state machine start
    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._StateMachine\: process (\Clock\) 
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State\: \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._States\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_0\;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.number\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.flag\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.result\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.dataIn.0\: std_logic_vector(31 downto 0);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.1\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.2\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.3\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.4\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.5\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.return.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.6\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Finished\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.return\ <= to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.SimpleMemory.ReadEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.SimpleMemory.WriteEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\ <= to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_0\;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.number\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.flag\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.result\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.1\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.2\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.3\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.4\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.return.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.5\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.return.1\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.6\ := to_unsigned(0, 32);
            else 
                case \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State\ is 
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Finished\ <= true;
                        else 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Finished\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_2\ => 
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.number\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.number.parameter.In\;
                        -- Begin SimpleMemory read.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.SimpleMemory.ReadEnable\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.SimpleMemory.ReadEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.dataIn.0\ := \DataIn\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.0\ := ConvertStdLogicVectorToUInt32(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.dataIn.0\) + to_unsigned(1, 32);
                            -- Begin SimpleMemory write.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.SimpleMemory.WriteEnable\ <= true;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.SimpleMemory.DataOut\ <= ConvertUInt32ToStdLogicVector(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.0\);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_4\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.SimpleMemory.WriteEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.1\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.number\ = to_signed(0, 16);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.2\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.number\ = to_signed(1, 16);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.3\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.1\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.2\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.flag\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.3\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_6\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_6\.
                            --     * The false branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_7\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_11\.
                            --     * Execution after either branch will continue in the following state: \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_5\.

                            if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.flag\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_6\;
                            else 
                                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_7\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_5\ => 
                        -- State after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.return\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.result\;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_6\ => 
                        -- True branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.result\ := resize(unsigned(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.number\), 32);
                        -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_4\.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_6\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_7\ => 
                        -- False branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.4\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.number\ - to_signed(2, 16);
                        -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.4\;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_8\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_8\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.return.0\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.5\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.number\ - to_signed(1, 16);
                            -- The last invocation for the target state machine just finished, so need to start the next one in a later state.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_9\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_9\ => 
                        -- This state was just added to leave time for the invocation proxy to register that the previous invocation finished.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_10\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_10\ => 
                        -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.5\;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_11\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_11\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.return.1\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.6\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.return.0\ + \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.return.1\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.result\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.binaryOperationResult.6\;
                            -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_4\.
                            if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_11\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._State_5\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).3 state machine end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).4 state machine start
    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._StateMachine\: process (\Clock\) 
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State\: \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._States\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_0\;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.number\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.flag\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.result\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.dataIn.0\: std_logic_vector(31 downto 0);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.1\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.2\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.3\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.4\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.5\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.return.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.6\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Finished\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.return\ <= to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.SimpleMemory.ReadEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.SimpleMemory.WriteEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\ <= to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_0\;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.number\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.flag\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.result\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.1\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.2\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.3\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.4\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.return.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.5\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.return.1\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.6\ := to_unsigned(0, 32);
            else 
                case \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State\ is 
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Finished\ <= true;
                        else 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Finished\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_2\ => 
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.number\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.number.parameter.In\;
                        -- Begin SimpleMemory read.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.SimpleMemory.ReadEnable\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.SimpleMemory.ReadEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.dataIn.0\ := \DataIn\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.0\ := ConvertStdLogicVectorToUInt32(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.dataIn.0\) + to_unsigned(1, 32);
                            -- Begin SimpleMemory write.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.SimpleMemory.WriteEnable\ <= true;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.SimpleMemory.DataOut\ <= ConvertUInt32ToStdLogicVector(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.0\);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_4\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.SimpleMemory.WriteEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.1\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.number\ = to_signed(0, 16);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.2\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.number\ = to_signed(1, 16);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.3\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.1\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.2\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.flag\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.3\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_6\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_6\.
                            --     * The false branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_7\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_11\.
                            --     * Execution after either branch will continue in the following state: \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_5\.

                            if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.flag\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_6\;
                            else 
                                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_7\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_5\ => 
                        -- State after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.return\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.result\;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_6\ => 
                        -- True branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.result\ := resize(unsigned(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.number\), 32);
                        -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_4\.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_6\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_7\ => 
                        -- False branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.4\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.number\ - to_signed(2, 16);
                        -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.4\;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_8\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_8\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.return.0\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.5\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.number\ - to_signed(1, 16);
                            -- The last invocation for the target state machine just finished, so need to start the next one in a later state.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_9\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_9\ => 
                        -- This state was just added to leave time for the invocation proxy to register that the previous invocation finished.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_10\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_10\ => 
                        -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.5\;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_11\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_11\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.return.1\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.6\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.return.0\ + \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.return.1\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.result\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.binaryOperationResult.6\;
                            -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_4\.
                            if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_11\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._State_5\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).4 state machine end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).5 state machine start
    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._StateMachine\: process (\Clock\) 
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State\: \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._States\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_0\;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.number\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.flag\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.result\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.dataIn.0\: std_logic_vector(31 downto 0);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.1\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.2\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.3\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.4\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.5\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.return.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.6\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Finished\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.return\ <= to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.SimpleMemory.ReadEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.SimpleMemory.WriteEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\ <= to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_0\;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.number\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.flag\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.result\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.1\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.2\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.3\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.4\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.return.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.5\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.return.1\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.6\ := to_unsigned(0, 32);
            else 
                case \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State\ is 
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Finished\ <= true;
                        else 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Finished\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_2\ => 
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.number\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.number.parameter.In\;
                        -- Begin SimpleMemory read.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.SimpleMemory.ReadEnable\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.SimpleMemory.ReadEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.dataIn.0\ := \DataIn\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.0\ := ConvertStdLogicVectorToUInt32(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.dataIn.0\) + to_unsigned(1, 32);
                            -- Begin SimpleMemory write.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.SimpleMemory.WriteEnable\ <= true;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.SimpleMemory.DataOut\ <= ConvertUInt32ToStdLogicVector(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.0\);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_4\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.SimpleMemory.WriteEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.1\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.number\ = to_signed(0, 16);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.2\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.number\ = to_signed(1, 16);
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.3\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.1\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.2\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.flag\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.3\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_6\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_6\.
                            --     * The false branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_7\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_11\.
                            --     * Execution after either branch will continue in the following state: \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_5\.

                            if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.flag\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_6\;
                            else 
                                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_7\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_5\ => 
                        -- State after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.return\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.result\;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_6\ => 
                        -- True branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.result\ := resize(unsigned(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.number\), 32);
                        -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_4\.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_6\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_7\ => 
                        -- False branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.4\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.number\ - to_signed(2, 16);
                        -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.4\;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_8\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_8\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.return.0\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.5\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.number\ - to_signed(1, 16);
                            -- The last invocation for the target state machine just finished, so need to start the next one in a later state.
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_9\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_9\ => 
                        -- This state was just added to leave time for the invocation proxy to register that the previous invocation finished.
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_10\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_10\ => 
                        -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.5\;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_11\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_11\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.return.1\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.6\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.return.0\ + \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.return.1\;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.result\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.binaryOperationResult.6\;
                            -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_4\.
                            if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State\ = \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_11\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._State_5\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).5 state machine end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).0 state machine start
    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._StateMachine\: process (\Clock\) 
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State\: \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._States\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_0\;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.number\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.flag\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.result\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.dataIn.0\: std_logic_vector(31 downto 0);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.binaryOperationResult.1\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.binaryOperationResult.2\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Finished\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.return\ <= to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.SimpleMemory.ReadEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.SimpleMemory.WriteEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\ <= to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_0\;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.number\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.flag\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.result\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.binaryOperationResult.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.binaryOperationResult.1\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.binaryOperationResult.2\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.return.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.binaryOperationResult.3\ := to_unsigned(0, 32);
            else 
                case \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State\ is 
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Finished\ <= true;
                        else 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Finished\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_2\ => 
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.number\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.number.parameter.In\;
                        -- Begin SimpleMemory read.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.SimpleMemory.ReadEnable\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.SimpleMemory.ReadEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.dataIn.0\ := \DataIn\;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.binaryOperationResult.0\ := ConvertStdLogicVectorToUInt32(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.dataIn.0\) + to_unsigned(1, 32);
                            -- Begin SimpleMemory write.
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.SimpleMemory.WriteEnable\ <= true;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.SimpleMemory.DataOut\ <= ConvertUInt32ToStdLogicVector(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.binaryOperationResult.0\);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_4\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.SimpleMemory.WriteEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.binaryOperationResult.1\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.number\ = to_signed(0, 16);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.flag\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.binaryOperationResult.1\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_6\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_6\.
                            --     * The false branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_7\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_8\.
                            --     * Execution after either branch will continue in the following state: \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_5\.

                            if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.flag\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_6\;
                            else 
                                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_7\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_5\ => 
                        -- State after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.return\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.result\;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_6\ => 
                        -- True branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.result\ := to_unsigned(1, 32);
                        -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_4\.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State\ = \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_6\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_7\ => 
                        -- False branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.binaryOperationResult.2\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.number\ - to_signed(1, 16);
                        -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.binaryOperationResult.2\;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_8\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_8\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ = \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.return.0\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.binaryOperationResult.3\ := resize(unsigned(resize(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.number\, 64) * signed((resize(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.return.0\, 64)))), 32);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.result\ := (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.binaryOperationResult.3\);
                            -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_4\.
                            if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State\ = \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_8\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._State_5\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).0 state machine end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).1 state machine start
    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._StateMachine\: process (\Clock\) 
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State\: \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._States\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_0\;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.number\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.flag\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.result\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.dataIn.0\: std_logic_vector(31 downto 0);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.binaryOperationResult.1\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.binaryOperationResult.2\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Finished\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.return\ <= to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.SimpleMemory.ReadEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.SimpleMemory.WriteEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\ <= to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_0\;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.number\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.flag\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.result\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.binaryOperationResult.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.binaryOperationResult.1\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.binaryOperationResult.2\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.return.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.binaryOperationResult.3\ := to_unsigned(0, 32);
            else 
                case \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State\ is 
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Finished\ <= true;
                        else 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Finished\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_2\ => 
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.number\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.number.parameter.In\;
                        -- Begin SimpleMemory read.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.SimpleMemory.ReadEnable\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.SimpleMemory.ReadEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.dataIn.0\ := \DataIn\;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.binaryOperationResult.0\ := ConvertStdLogicVectorToUInt32(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.dataIn.0\) + to_unsigned(1, 32);
                            -- Begin SimpleMemory write.
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.SimpleMemory.WriteEnable\ <= true;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.SimpleMemory.DataOut\ <= ConvertUInt32ToStdLogicVector(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.binaryOperationResult.0\);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_4\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.SimpleMemory.WriteEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.binaryOperationResult.1\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.number\ = to_signed(0, 16);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.flag\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.binaryOperationResult.1\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_6\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_6\.
                            --     * The false branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_7\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_8\.
                            --     * Execution after either branch will continue in the following state: \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_5\.

                            if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.flag\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_6\;
                            else 
                                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_7\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_5\ => 
                        -- State after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.return\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.result\;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_6\ => 
                        -- True branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.result\ := to_unsigned(1, 32);
                        -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_4\.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State\ = \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_6\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_7\ => 
                        -- False branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.binaryOperationResult.2\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.number\ - to_signed(1, 16);
                        -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.binaryOperationResult.2\;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_8\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_8\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ = \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.return.0\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.binaryOperationResult.3\ := resize(unsigned(resize(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.number\, 64) * signed((resize(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.return.0\, 64)))), 32);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.result\ := (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.binaryOperationResult.3\);
                            -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_4\.
                            if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State\ = \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_8\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._State_5\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).1 state machine end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).2 state machine start
    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._StateMachine\: process (\Clock\) 
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State\: \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._States\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_0\;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.number\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.flag\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.result\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.dataIn.0\: std_logic_vector(31 downto 0);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.binaryOperationResult.1\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.binaryOperationResult.2\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Finished\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.return\ <= to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.SimpleMemory.ReadEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.SimpleMemory.WriteEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\ <= to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_0\;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.number\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.flag\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.result\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.binaryOperationResult.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.binaryOperationResult.1\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.binaryOperationResult.2\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.return.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.binaryOperationResult.3\ := to_unsigned(0, 32);
            else 
                case \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State\ is 
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Finished\ <= true;
                        else 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Finished\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_2\ => 
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.number\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.number.parameter.In\;
                        -- Begin SimpleMemory read.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.SimpleMemory.ReadEnable\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.SimpleMemory.ReadEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.dataIn.0\ := \DataIn\;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.binaryOperationResult.0\ := ConvertStdLogicVectorToUInt32(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.dataIn.0\) + to_unsigned(1, 32);
                            -- Begin SimpleMemory write.
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.SimpleMemory.WriteEnable\ <= true;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.SimpleMemory.DataOut\ <= ConvertUInt32ToStdLogicVector(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.binaryOperationResult.0\);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_4\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.SimpleMemory.WriteEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.binaryOperationResult.1\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.number\ = to_signed(0, 16);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.flag\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.binaryOperationResult.1\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_6\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_6\.
                            --     * The false branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_7\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_8\.
                            --     * Execution after either branch will continue in the following state: \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_5\.

                            if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.flag\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_6\;
                            else 
                                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_7\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_5\ => 
                        -- State after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.return\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.result\;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_6\ => 
                        -- True branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.result\ := to_unsigned(1, 32);
                        -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_4\.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State\ = \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_6\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_7\ => 
                        -- False branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.binaryOperationResult.2\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.number\ - to_signed(1, 16);
                        -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.binaryOperationResult.2\;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_8\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_8\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ = \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.return.0\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.binaryOperationResult.3\ := resize(unsigned(resize(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.number\, 64) * signed((resize(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.return.0\, 64)))), 32);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.result\ := (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.binaryOperationResult.3\);
                            -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_4\.
                            if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State\ = \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_8\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._State_5\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).2 state machine end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).3 state machine start
    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._StateMachine\: process (\Clock\) 
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State\: \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._States\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_0\;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.number\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.flag\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.result\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.dataIn.0\: std_logic_vector(31 downto 0);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.binaryOperationResult.1\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.binaryOperationResult.2\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Finished\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.return\ <= to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.SimpleMemory.ReadEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.SimpleMemory.WriteEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\ <= to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_0\;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.number\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.flag\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.result\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.binaryOperationResult.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.binaryOperationResult.1\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.binaryOperationResult.2\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.return.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.binaryOperationResult.3\ := to_unsigned(0, 32);
            else 
                case \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State\ is 
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Finished\ <= true;
                        else 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Finished\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_2\ => 
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.number\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.number.parameter.In\;
                        -- Begin SimpleMemory read.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.SimpleMemory.ReadEnable\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.SimpleMemory.ReadEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.dataIn.0\ := \DataIn\;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.binaryOperationResult.0\ := ConvertStdLogicVectorToUInt32(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.dataIn.0\) + to_unsigned(1, 32);
                            -- Begin SimpleMemory write.
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.SimpleMemory.WriteEnable\ <= true;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.SimpleMemory.DataOut\ <= ConvertUInt32ToStdLogicVector(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.binaryOperationResult.0\);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_4\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.SimpleMemory.WriteEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.binaryOperationResult.1\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.number\ = to_signed(0, 16);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.flag\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.binaryOperationResult.1\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_6\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_6\.
                            --     * The false branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_7\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_8\.
                            --     * Execution after either branch will continue in the following state: \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_5\.

                            if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.flag\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_6\;
                            else 
                                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_7\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_5\ => 
                        -- State after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.return\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.result\;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_6\ => 
                        -- True branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.result\ := to_unsigned(1, 32);
                        -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_4\.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State\ = \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_6\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_7\ => 
                        -- False branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.binaryOperationResult.2\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.number\ - to_signed(1, 16);
                        -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.binaryOperationResult.2\;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_8\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_8\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ = \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.return.0\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.binaryOperationResult.3\ := resize(unsigned(resize(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.number\, 64) * signed((resize(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.return.0\, 64)))), 32);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.result\ := (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.binaryOperationResult.3\);
                            -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_4\.
                            if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State\ = \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_8\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._State_5\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).3 state machine end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).4 state machine start
    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._StateMachine\: process (\Clock\) 
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State\: \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._States\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_0\;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.number\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.flag\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.result\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.dataIn.0\: std_logic_vector(31 downto 0);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.binaryOperationResult.1\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.binaryOperationResult.2\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Finished\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.return\ <= to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.SimpleMemory.ReadEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.SimpleMemory.WriteEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\ <= to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_0\;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.number\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.flag\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.result\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.binaryOperationResult.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.binaryOperationResult.1\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.binaryOperationResult.2\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.return.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.binaryOperationResult.3\ := to_unsigned(0, 32);
            else 
                case \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State\ is 
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Finished\ <= true;
                        else 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Finished\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_2\ => 
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.number\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.number.parameter.In\;
                        -- Begin SimpleMemory read.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.SimpleMemory.ReadEnable\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.SimpleMemory.ReadEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.dataIn.0\ := \DataIn\;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.binaryOperationResult.0\ := ConvertStdLogicVectorToUInt32(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.dataIn.0\) + to_unsigned(1, 32);
                            -- Begin SimpleMemory write.
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.SimpleMemory.WriteEnable\ <= true;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.SimpleMemory.DataOut\ <= ConvertUInt32ToStdLogicVector(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.binaryOperationResult.0\);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_4\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.SimpleMemory.WriteEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.binaryOperationResult.1\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.number\ = to_signed(0, 16);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.flag\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.binaryOperationResult.1\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_6\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_6\.
                            --     * The false branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_7\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_8\.
                            --     * Execution after either branch will continue in the following state: \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_5\.

                            if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.flag\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_6\;
                            else 
                                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_7\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_5\ => 
                        -- State after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.return\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.result\;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_6\ => 
                        -- True branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.result\ := to_unsigned(1, 32);
                        -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_4\.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State\ = \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_6\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_7\ => 
                        -- False branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.binaryOperationResult.2\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.number\ - to_signed(1, 16);
                        -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.binaryOperationResult.2\;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_8\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_8\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ = \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.return.0\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.binaryOperationResult.3\ := resize(unsigned(resize(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.number\, 64) * signed((resize(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.return.0\, 64)))), 32);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.result\ := (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.binaryOperationResult.3\);
                            -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_4\.
                            if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State\ = \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_8\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._State_5\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).4 state machine end


    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).5 state machine start
    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._StateMachine\: process (\Clock\) 
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State\: \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._States\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_0\;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.number\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.flag\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.result\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.dataIn.0\: std_logic_vector(31 downto 0);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.binaryOperationResult.1\: boolean := false;
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.binaryOperationResult.2\: signed(15 downto 0) := to_signed(0, 16);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Finished\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.return\ <= to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.SimpleMemory.ReadEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.SimpleMemory.WriteEnable\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\ <= to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_0\;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.number\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.flag\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.result\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.binaryOperationResult.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.binaryOperationResult.1\ := false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.binaryOperationResult.2\ := to_signed(0, 16);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.return.0\ := to_unsigned(0, 32);
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.binaryOperationResult.3\ := to_unsigned(0, 32);
            else 
                case \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State\ is 
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Started\ = true) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Finished\ <= true;
                        else 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Finished\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_2\ => 
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.number\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.number.parameter.In\;
                        -- Begin SimpleMemory read.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.SimpleMemory.ReadEnable\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.SimpleMemory.ReadEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.dataIn.0\ := \DataIn\;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.binaryOperationResult.0\ := ConvertStdLogicVectorToUInt32(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.dataIn.0\) + to_unsigned(1, 32);
                            -- Begin SimpleMemory write.
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.SimpleMemory.CellIndex\ <= resize(to_signed(1, 32), 32);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.SimpleMemory.WriteEnable\ <= true;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.SimpleMemory.DataOut\ <= ConvertUInt32ToStdLogicVector(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.binaryOperationResult.0\);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_4\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.SimpleMemory.WriteEnable\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.binaryOperationResult.1\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.number\ = to_signed(0, 16);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.flag\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.binaryOperationResult.1\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_6\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_6\.
                            --     * The false branch starts in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_7\ and ends in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_8\.
                            --     * Execution after either branch will continue in the following state: \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_5\.

                            if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.flag\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_6\;
                            else 
                                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_7\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_5\ => 
                        -- State after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.return\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.result\;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_6\ => 
                        -- True branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.result\ := to_unsigned(1, 32);
                        -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_4\.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State\ = \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_6\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_7\ => 
                        -- False branch of the if-else started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_4\.
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.binaryOperationResult.2\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.number\ - to_signed(1, 16);
                        -- Starting state machine invocation for the following method: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.binaryOperationResult.2\;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ <= true;
                        \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_8\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_8\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16)
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ = \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ <= false;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.return.0\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.binaryOperationResult.3\ := resize(unsigned(resize(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.number\, 64) * signed((resize(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.return.0\, 64)))), 32);
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.result\ := (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.binaryOperationResult.3\);
                            -- Going to the state after the if-else which was started in state \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_4\.
                            if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State\ = \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_8\) then 
                                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State\ := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._State_5\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).5 state machine end


    -- System.Void Hast.Samples.SampleAssembly.SimdCalculator::AddVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine start
    \SimdCalculator::AddVectors(SimpleMemory).0._StateMachine\: process (\Clock\) 
        Variable \SimdCalculator::AddVectors(SimpleMemory).0._State\: \SimdCalculator::AddVectors(SimpleMemory).0._States\ := \SimdCalculator::AddVectors(SimpleMemory).0._State_0\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \SimdCalculator::AddVectors(SimpleMemory).0._Finished\ <= false;
                \SimdCalculator::AddVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\ <= false;
                \SimdCalculator::AddVectors(SimpleMemory).0._State\ := \SimdCalculator::AddVectors(SimpleMemory).0._State_0\;
            else 
                case \SimdCalculator::AddVectors(SimpleMemory).0._State\ is 
                    when \SimdCalculator::AddVectors(SimpleMemory).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\SimdCalculator::AddVectors(SimpleMemory).0._Started\ = true) then 
                            \SimdCalculator::AddVectors(SimpleMemory).0._State\ := \SimdCalculator::AddVectors(SimpleMemory).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \SimdCalculator::AddVectors(SimpleMemory).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\SimdCalculator::AddVectors(SimpleMemory).0._Started\ = true) then 
                            \SimdCalculator::AddVectors(SimpleMemory).0._Finished\ <= true;
                        else 
                            \SimdCalculator::AddVectors(SimpleMemory).0._Finished\ <= false;
                            \SimdCalculator::AddVectors(SimpleMemory).0._State\ := \SimdCalculator::AddVectors(SimpleMemory).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \SimdCalculator::AddVectors(SimpleMemory).0._State_2\ => 
                        -- Starting state machine invocation for the following method: System.Void Hast.Samples.SampleAssembly.SimdCalculator::RunSimdOperation(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,Hast.Samples.SampleAssembly.SimdOperation)
                        \SimdCalculator::AddVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).operation.parameter.Out.0\ <= \Hast.Samples.SampleAssembly.SimdOperation Hast.Samples.SampleAssembly.SimdOperation::Add\;
                        \SimdCalculator::AddVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\ <= true;
                        \SimdCalculator::AddVectors(SimpleMemory).0._State\ := \SimdCalculator::AddVectors(SimpleMemory).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \SimdCalculator::AddVectors(SimpleMemory).0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.Samples.SampleAssembly.SimdCalculator::RunSimdOperation(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,Hast.Samples.SampleAssembly.SimdOperation)
                        if (\SimdCalculator::AddVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\ = \SimdCalculator::AddVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\) then 
                            \SimdCalculator::AddVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\ <= false;
                            \SimdCalculator::AddVectors(SimpleMemory).0._State\ := \SimdCalculator::AddVectors(SimpleMemory).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.Samples.SampleAssembly.SimdCalculator::AddVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine end


    -- System.Void Hast.Samples.SampleAssembly.SimdCalculator::SubtractVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine start
    \SimdCalculator::SubtractVectors(SimpleMemory).0._StateMachine\: process (\Clock\) 
        Variable \SimdCalculator::SubtractVectors(SimpleMemory).0._State\: \SimdCalculator::SubtractVectors(SimpleMemory).0._States\ := \SimdCalculator::SubtractVectors(SimpleMemory).0._State_0\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \SimdCalculator::SubtractVectors(SimpleMemory).0._Finished\ <= false;
                \SimdCalculator::SubtractVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\ <= false;
                \SimdCalculator::SubtractVectors(SimpleMemory).0._State\ := \SimdCalculator::SubtractVectors(SimpleMemory).0._State_0\;
            else 
                case \SimdCalculator::SubtractVectors(SimpleMemory).0._State\ is 
                    when \SimdCalculator::SubtractVectors(SimpleMemory).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\SimdCalculator::SubtractVectors(SimpleMemory).0._Started\ = true) then 
                            \SimdCalculator::SubtractVectors(SimpleMemory).0._State\ := \SimdCalculator::SubtractVectors(SimpleMemory).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \SimdCalculator::SubtractVectors(SimpleMemory).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\SimdCalculator::SubtractVectors(SimpleMemory).0._Started\ = true) then 
                            \SimdCalculator::SubtractVectors(SimpleMemory).0._Finished\ <= true;
                        else 
                            \SimdCalculator::SubtractVectors(SimpleMemory).0._Finished\ <= false;
                            \SimdCalculator::SubtractVectors(SimpleMemory).0._State\ := \SimdCalculator::SubtractVectors(SimpleMemory).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \SimdCalculator::SubtractVectors(SimpleMemory).0._State_2\ => 
                        -- Starting state machine invocation for the following method: System.Void Hast.Samples.SampleAssembly.SimdCalculator::RunSimdOperation(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,Hast.Samples.SampleAssembly.SimdOperation)
                        \SimdCalculator::SubtractVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).operation.parameter.Out.0\ <= \Hast.Samples.SampleAssembly.SimdOperation Hast.Samples.SampleAssembly.SimdOperation::Subtract\;
                        \SimdCalculator::SubtractVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\ <= true;
                        \SimdCalculator::SubtractVectors(SimpleMemory).0._State\ := \SimdCalculator::SubtractVectors(SimpleMemory).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \SimdCalculator::SubtractVectors(SimpleMemory).0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.Samples.SampleAssembly.SimdCalculator::RunSimdOperation(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,Hast.Samples.SampleAssembly.SimdOperation)
                        if (\SimdCalculator::SubtractVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\ = \SimdCalculator::SubtractVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\) then 
                            \SimdCalculator::SubtractVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\ <= false;
                            \SimdCalculator::SubtractVectors(SimpleMemory).0._State\ := \SimdCalculator::SubtractVectors(SimpleMemory).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.Samples.SampleAssembly.SimdCalculator::SubtractVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine end


    -- System.Void Hast.Samples.SampleAssembly.SimdCalculator::MultiplyVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine start
    \SimdCalculator::MultiplyVectors(SimpleMemory).0._StateMachine\: process (\Clock\) 
        Variable \SimdCalculator::MultiplyVectors(SimpleMemory).0._State\: \SimdCalculator::MultiplyVectors(SimpleMemory).0._States\ := \SimdCalculator::MultiplyVectors(SimpleMemory).0._State_0\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \SimdCalculator::MultiplyVectors(SimpleMemory).0._Finished\ <= false;
                \SimdCalculator::MultiplyVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\ <= false;
                \SimdCalculator::MultiplyVectors(SimpleMemory).0._State\ := \SimdCalculator::MultiplyVectors(SimpleMemory).0._State_0\;
            else 
                case \SimdCalculator::MultiplyVectors(SimpleMemory).0._State\ is 
                    when \SimdCalculator::MultiplyVectors(SimpleMemory).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\SimdCalculator::MultiplyVectors(SimpleMemory).0._Started\ = true) then 
                            \SimdCalculator::MultiplyVectors(SimpleMemory).0._State\ := \SimdCalculator::MultiplyVectors(SimpleMemory).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \SimdCalculator::MultiplyVectors(SimpleMemory).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\SimdCalculator::MultiplyVectors(SimpleMemory).0._Started\ = true) then 
                            \SimdCalculator::MultiplyVectors(SimpleMemory).0._Finished\ <= true;
                        else 
                            \SimdCalculator::MultiplyVectors(SimpleMemory).0._Finished\ <= false;
                            \SimdCalculator::MultiplyVectors(SimpleMemory).0._State\ := \SimdCalculator::MultiplyVectors(SimpleMemory).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \SimdCalculator::MultiplyVectors(SimpleMemory).0._State_2\ => 
                        -- Starting state machine invocation for the following method: System.Void Hast.Samples.SampleAssembly.SimdCalculator::RunSimdOperation(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,Hast.Samples.SampleAssembly.SimdOperation)
                        \SimdCalculator::MultiplyVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).operation.parameter.Out.0\ <= \Hast.Samples.SampleAssembly.SimdOperation Hast.Samples.SampleAssembly.SimdOperation::Multiply\;
                        \SimdCalculator::MultiplyVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\ <= true;
                        \SimdCalculator::MultiplyVectors(SimpleMemory).0._State\ := \SimdCalculator::MultiplyVectors(SimpleMemory).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \SimdCalculator::MultiplyVectors(SimpleMemory).0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.Samples.SampleAssembly.SimdCalculator::RunSimdOperation(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,Hast.Samples.SampleAssembly.SimdOperation)
                        if (\SimdCalculator::MultiplyVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\ = \SimdCalculator::MultiplyVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\) then 
                            \SimdCalculator::MultiplyVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\ <= false;
                            \SimdCalculator::MultiplyVectors(SimpleMemory).0._State\ := \SimdCalculator::MultiplyVectors(SimpleMemory).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.Samples.SampleAssembly.SimdCalculator::MultiplyVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine end


    -- System.Void Hast.Samples.SampleAssembly.SimdCalculator::DivideVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine start
    \SimdCalculator::DivideVectors(SimpleMemory).0._StateMachine\: process (\Clock\) 
        Variable \SimdCalculator::DivideVectors(SimpleMemory).0._State\: \SimdCalculator::DivideVectors(SimpleMemory).0._States\ := \SimdCalculator::DivideVectors(SimpleMemory).0._State_0\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \SimdCalculator::DivideVectors(SimpleMemory).0._Finished\ <= false;
                \SimdCalculator::DivideVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\ <= false;
                \SimdCalculator::DivideVectors(SimpleMemory).0._State\ := \SimdCalculator::DivideVectors(SimpleMemory).0._State_0\;
            else 
                case \SimdCalculator::DivideVectors(SimpleMemory).0._State\ is 
                    when \SimdCalculator::DivideVectors(SimpleMemory).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\SimdCalculator::DivideVectors(SimpleMemory).0._Started\ = true) then 
                            \SimdCalculator::DivideVectors(SimpleMemory).0._State\ := \SimdCalculator::DivideVectors(SimpleMemory).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \SimdCalculator::DivideVectors(SimpleMemory).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\SimdCalculator::DivideVectors(SimpleMemory).0._Started\ = true) then 
                            \SimdCalculator::DivideVectors(SimpleMemory).0._Finished\ <= true;
                        else 
                            \SimdCalculator::DivideVectors(SimpleMemory).0._Finished\ <= false;
                            \SimdCalculator::DivideVectors(SimpleMemory).0._State\ := \SimdCalculator::DivideVectors(SimpleMemory).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \SimdCalculator::DivideVectors(SimpleMemory).0._State_2\ => 
                        -- Starting state machine invocation for the following method: System.Void Hast.Samples.SampleAssembly.SimdCalculator::RunSimdOperation(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,Hast.Samples.SampleAssembly.SimdOperation)
                        \SimdCalculator::DivideVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).operation.parameter.Out.0\ <= \Hast.Samples.SampleAssembly.SimdOperation Hast.Samples.SampleAssembly.SimdOperation::Divide\;
                        \SimdCalculator::DivideVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\ <= true;
                        \SimdCalculator::DivideVectors(SimpleMemory).0._State\ := \SimdCalculator::DivideVectors(SimpleMemory).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \SimdCalculator::DivideVectors(SimpleMemory).0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.Samples.SampleAssembly.SimdCalculator::RunSimdOperation(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,Hast.Samples.SampleAssembly.SimdOperation)
                        if (\SimdCalculator::DivideVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\ = \SimdCalculator::DivideVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\) then 
                            \SimdCalculator::DivideVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\ <= false;
                            \SimdCalculator::DivideVectors(SimpleMemory).0._State\ := \SimdCalculator::DivideVectors(SimpleMemory).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.Samples.SampleAssembly.SimdCalculator::DivideVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine end


    -- System.Void Hast.Samples.SampleAssembly.SimdCalculator::RunSimdOperation(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,Hast.Samples.SampleAssembly.SimdOperation).0 state machine start
    \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._StateMachine\: process (\Clock\) 
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\: \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._States\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_0\;
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.operation\: \Hast.Samples.SampleAssembly.SimdOperation\;
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.num\: signed(31 downto 0) := to_signed(0, 32);
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.i\: signed(31 downto 0) := to_signed(0, 32);
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\: \signed32_Array\(0 to 29) := (others => to_signed(0, 32));
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\: \signed32_Array\(0 to 29) := (others => to_signed(0, 32));
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array3\: \signed32_Array\(0 to 29) := (others => to_signed(0, 32));
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.j\: signed(31 downto 0) := to_signed(0, 32);
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.k\: signed(31 downto 0) := to_signed(0, 32);
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.l\: signed(31 downto 0) := to_signed(0, 32);
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.dataIn.0\: std_logic_vector(31 downto 0);
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.0\: boolean := false;
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.1\: boolean := false;
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.2\: boolean := false;
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.3\: boolean := false;
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.4\: signed(31 downto 0) := to_signed(0, 32);
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.5\: signed(31 downto 0) := to_signed(0, 32);
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.dataIn.1\: std_logic_vector(31 downto 0);
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.6\: signed(31 downto 0) := to_signed(0, 32);
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.7\: boolean := false;
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.8\: boolean := false;
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.9\: signed(31 downto 0) := to_signed(0, 32);
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.10\: signed(31 downto 0) := to_signed(0, 32);
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.11\: signed(31 downto 0) := to_signed(0, 32);
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.dataIn.2\: std_logic_vector(31 downto 0);
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.12\: signed(31 downto 0) := to_signed(0, 32);
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.133\: boolean := false;
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.134\: boolean := false;
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.135\: signed(31 downto 0) := to_signed(0, 32);
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.136\: signed(31 downto 0) := to_signed(0, 32);
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.137\: signed(31 downto 0) := to_signed(0, 32);
        Variable \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.138\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._Finished\ <= false;
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.ReadEnable\ <= false;
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.WriteEnable\ <= false;
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.13\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.14\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.15\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.16\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.17\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.18\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.19\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.20\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.21\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.22\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.23\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.24\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.25\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.26\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.27\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.28\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.29\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.30\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.31\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.32\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.33\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.34\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.35\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.36\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.37\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.38\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.39\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.40\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.41\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.42\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.43\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.44\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.45\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.46\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.47\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.48\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.49\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.50\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.51\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.52\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.53\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.54\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.55\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.56\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.57\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.58\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.59\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.60\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.61\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.62\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.63\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.64\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.65\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.66\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.67\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.68\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.69\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.70\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.71\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.72\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.73\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.74\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.75\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.76\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.77\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.78\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.79\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.80\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.81\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.82\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.83\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.84\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.85\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.86\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.87\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.88\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.89\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.90\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.91\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.92\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.93\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.94\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.95\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.96\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.97\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.98\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.99\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.100\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.101\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.102\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.103\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.104\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.105\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.106\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.107\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.108\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.109\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.110\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.111\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.112\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.113\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.114\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.115\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.116\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.117\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.118\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.119\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.120\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.121\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.122\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.123\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.124\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.125\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.126\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.127\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.128\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.129\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.130\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.131\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.132\ <= to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_0\;
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.num\ := to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.i\ := to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\ := (others => to_signed(0, 32));
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\ := (others => to_signed(0, 32));
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array3\ := (others => to_signed(0, 32));
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.j\ := to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.k\ := to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.l\ := to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.0\ := false;
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.1\ := false;
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.2\ := false;
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.3\ := false;
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.4\ := to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.5\ := to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.6\ := to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.7\ := false;
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.8\ := false;
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.9\ := to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.10\ := to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.11\ := to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.12\ := to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.133\ := false;
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.134\ := false;
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.135\ := to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.136\ := to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.137\ := to_signed(0, 32);
                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.138\ := to_signed(0, 32);
            else 
                case \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ is 
                    when \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._Started\ = true) then 
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._Started\ = true) then 
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._Finished\ <= true;
                        else 
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._Finished\ <= false;
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_2\ => 
                        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.operation\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.operation.parameter.In\;
                        -- Begin SimpleMemory read.
                        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.CellIndex\ <= resize(to_signed(0, 32), 32);
                        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.ReadEnable\ <= true;
                        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.ReadEnable\ <= false;
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.dataIn.0\ := \DataIn\;
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.num\ := ConvertStdLogicVectorToInt32(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.dataIn.0\);
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.i\ := to_signed(0, 32);
                            -- Starting a while loop.
                            -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.0\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.i\ < \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.num\;
                            if (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.0\) then 
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_4\;
                            else 
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_5\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_4\ => 
                        -- Repeated state of the while loop which was started in state \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_3\.
                        -- The while loop's condition:
                        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.1\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.i\ < \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.num\;
                        if (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.1\) then 
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\ := (others => to_signed(0, 32));
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\ := (others => to_signed(0, 32));
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array3\ := (others => to_signed(0, 32));
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.j\ := to_signed(0, 32);
                            -- Starting a while loop.
                            -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.2\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.j\ < to_signed(30, 32);
                            if (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.2\) then 
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_6\;
                            else 
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_7\;
                            end if;
                        else 
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_5\ => 
                        -- State after the while loop which was started in state \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_3\.
                        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_6\ => 
                        -- Repeated state of the while loop which was started in state \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_4\.
                        -- The while loop's condition:
                        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.3\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.j\ < to_signed(30, 32);
                        if (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.3\) then 
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.4\ := to_signed(1, 32) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.i\;
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.5\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.4\ + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.j\;
                            -- Begin SimpleMemory read.
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.CellIndex\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.5\, 32);
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.ReadEnable\ <= true;
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_8\;
                        else 
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_7\ => 
                        -- State after the while loop which was started in state \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_4\.
                        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.k\ := to_signed(0, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.7\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.k\ < to_signed(30, 32);
                        if (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.7\) then 
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_9\;
                        else 
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_10\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_8\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.ReadEnable\ <= false;
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.dataIn.1\ := \DataIn\;
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(to_integer(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.j\)) := ConvertStdLogicVectorToInt32(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.dataIn.1\);
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.6\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.j\ + to_signed(1, 32);
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.j\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.6\;
                            -- Returning to the repeated state of the while loop which was started in state \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_4\ if the loop wasn't exited with a state change.
                            if (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ = \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_8\) then 
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_6\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_9\ => 
                        -- Repeated state of the while loop which was started in state \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_7\.
                        -- The while loop's condition:
                        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.8\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.k\ < to_signed(30, 32);
                        if (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.8\) then 
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.9\ := to_signed(1, 32) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.i\;
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.10\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.9\ + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.k\;
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.11\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.10\ + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.num\;
                            -- Begin SimpleMemory read.
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.CellIndex\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.11\, 32);
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.ReadEnable\ <= true;
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_11\;
                        else 
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_10\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.4
                    when \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_10\ => 
                        -- State after the while loop which was started in state \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_7\.
                        case \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.operation\ is 
                            when \Hast.Samples.SampleAssembly.SimdOperation Hast.Samples.SampleAssembly.SimdOperation::Add\ => 
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.13\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(0) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(0);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.14\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(1) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(1);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.15\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(2) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(2);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.16\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(3) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(3);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.17\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(4) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(4);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.18\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(5) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(5);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.19\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(6) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(6);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.20\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(7) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(7);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.21\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(8) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(8);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.22\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(9) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(9);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.23\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(10) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(10);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.24\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(11) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(11);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.25\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(12) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(12);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.26\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(13) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(13);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.27\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(14) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(14);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.28\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(15) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(15);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.29\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(16) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(16);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.30\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(17) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(17);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.31\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(18) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(18);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.32\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(19) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(19);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.33\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(20) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(20);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.34\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(21) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(21);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.35\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(22) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(22);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.36\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(23) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(23);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.37\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(24) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(24);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.38\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(25) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(25);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.39\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(26) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(26);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.40\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(27) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(27);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.41\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(28) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(28);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.42\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(29) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(29);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_13\;
                            when \Hast.Samples.SampleAssembly.SimdOperation Hast.Samples.SampleAssembly.SimdOperation::Subtract\ => 
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.43\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(0) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(0);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.44\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(1) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(1);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.45\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(2) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(2);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.46\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(3) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(3);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.47\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(4) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(4);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.48\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(5) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(5);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.49\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(6) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(6);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.50\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(7) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(7);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.51\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(8) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(8);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.52\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(9) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(9);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.53\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(10) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(10);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.54\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(11) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(11);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.55\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(12) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(12);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.56\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(13) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(13);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.57\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(14) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(14);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.58\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(15) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(15);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.59\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(16) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(16);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.60\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(17) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(17);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.61\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(18) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(18);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.62\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(19) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(19);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.63\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(20) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(20);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.64\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(21) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(21);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.65\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(22) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(22);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.66\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(23) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(23);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.67\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(24) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(24);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.68\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(25) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(25);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.69\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(26) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(26);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.70\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(27) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(27);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.71\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(28) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(28);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.72\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(29) - \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(29);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_14\;
                            when \Hast.Samples.SampleAssembly.SimdOperation Hast.Samples.SampleAssembly.SimdOperation::Multiply\ => 
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.73\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(0) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(0), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.74\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(1) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(1), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.75\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(2) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(2), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.76\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(3) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(3), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.77\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(4) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(4), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.78\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(5) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(5), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.79\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(6) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(6), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.80\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(7) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(7), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.81\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(8) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(8), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.82\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(9) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(9), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.83\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(10) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(10), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.84\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(11) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(11), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.85\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(12) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(12), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.86\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(13) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(13), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.87\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(14) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(14), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.88\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(15) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(15), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.89\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(16) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(16), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.90\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(17) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(17), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.91\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(18) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(18), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.92\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(19) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(19), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.93\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(20) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(20), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.94\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(21) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(21), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.95\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(22) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(22), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.96\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(23) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(23), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.97\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(24) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(24), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.98\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(25) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(25), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.99\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(26) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(26), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.100\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(27) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(27), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.101\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(28) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(28), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.102\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(29) * \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(29), 32);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_15\;
                            when \Hast.Samples.SampleAssembly.SimdOperation Hast.Samples.SampleAssembly.SimdOperation::Divide\ => 
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.103\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(0) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(0);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.104\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(1) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(1);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.105\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(2) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(2);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.106\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(3) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(3);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.107\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(4) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(4);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.108\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(5) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(5);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.109\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(6) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(6);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.110\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(7) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(7);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.111\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(8) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(8);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.112\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(9) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(9);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.113\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(10) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(10);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.114\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(11) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(11);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.115\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(12) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(12);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.116\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(13) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(13);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.117\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(14) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(14);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.118\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(15) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(15);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.119\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(16) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(16);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.120\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(17) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(17);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.121\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(18) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(18);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.122\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(19) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(19);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.123\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(20) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(20);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.124\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(21) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(21);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.125\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(22) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(22);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.126\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(23) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(23);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.127\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(24) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(24);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.128\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(25) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(25);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.129\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(26) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(26);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.130\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(27) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(27);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.131\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(28) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(28);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.132\ <= \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array\(29) / \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(29);
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_16\;
                        end case;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_11\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.ReadEnable\ <= false;
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.dataIn.2\ := \DataIn\;
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array2\(to_integer(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.k\)) := ConvertStdLogicVectorToInt32(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.dataIn.2\);
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.12\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.k\ + to_signed(1, 32);
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.k\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.12\;
                            -- Returning to the repeated state of the while loop which was started in state \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_7\ if the loop wasn't exited with a state change.
                            if (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ = \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_11\) then 
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_9\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_12\ => 
                        -- State after the case statement which was started in state \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_10\.
                        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.l\ := to_signed(0, 32);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.133\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.l\ < to_signed(30, 32);
                        if (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.133\) then 
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_17\;
                        else 
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_18\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_13\ => 
                        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array3\ := (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.13\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.14\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.15\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.16\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.17\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.18\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.19\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.20\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.21\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.22\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.23\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.24\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.25\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.26\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.27\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.28\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.29\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.30\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.31\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.32\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.33\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.34\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.35\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.36\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.37\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.38\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.39\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.40\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.41\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.42\);
                        -- Going to the state after the case statement which was started in state \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_10\.
                        if (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ = \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_13\) then 
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_12\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_14\ => 
                        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array3\ := (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.43\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.44\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.45\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.46\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.47\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.48\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.49\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.50\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.51\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.52\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.53\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.54\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.55\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.56\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.57\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.58\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.59\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.60\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.61\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.62\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.63\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.64\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.65\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.66\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.67\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.68\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.69\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.70\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.71\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.72\);
                        -- Going to the state after the case statement which was started in state \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_10\.
                        if (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ = \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_14\) then 
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_12\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_15\ => 
                        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array3\ := (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.73\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.74\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.75\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.76\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.77\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.78\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.79\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.80\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.81\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.82\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.83\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.84\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.85\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.86\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.87\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.88\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.89\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.90\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.91\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.92\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.93\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.94\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.95\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.96\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.97\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.98\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.99\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.100\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.101\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.102\);
                        -- Going to the state after the case statement which was started in state \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_10\.
                        if (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ = \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_15\) then 
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_12\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_16\ => 
                        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array3\ := (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.103\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.104\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.105\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.106\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.107\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.108\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.109\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.110\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.111\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.112\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.113\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.114\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.115\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.116\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.117\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.118\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.119\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.120\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.121\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.122\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.123\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.124\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.125\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.126\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.127\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.128\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.129\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.130\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.131\, \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.132\);
                        -- Going to the state after the case statement which was started in state \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_10\.
                        if (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ = \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_16\) then 
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_12\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_17\ => 
                        -- Repeated state of the while loop which was started in state \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_12\.
                        -- The while loop's condition:
                        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.134\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.l\ < to_signed(30, 32);
                        if (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.134\) then 
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.135\ := to_signed(1, 32) + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.i\;
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.136\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.135\ + \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.l\;
                            -- Begin SimpleMemory write.
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.CellIndex\ <= resize(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.136\, 32);
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.WriteEnable\ <= true;
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.DataOut\ <= ConvertInt32ToStdLogicVector(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.array3\(to_integer(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.l\)));
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_19\;
                        else 
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_18\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_18\ => 
                        -- State after the while loop which was started in state \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_12\.
                        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.138\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.i\ + to_signed(30, 32);
                        \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.i\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.138\;
                        -- Returning to the repeated state of the while loop which was started in state \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_3\ if the loop wasn't exited with a state change.
                        if (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ = \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_18\) then 
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_19\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.WriteEnable\ <= false;
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.137\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.l\ + to_signed(1, 32);
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.l\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.binaryOperationResult.137\;
                            -- Returning to the repeated state of the while loop which was started in state \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_12\ if the loop wasn't exited with a state change.
                            if (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ = \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_19\) then 
                                \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State\ := \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._State_17\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.Samples.SampleAssembly.SimdCalculator::RunSimdOperation(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,Hast.Samples.SampleAssembly.SimdOperation).0 state machine end


    -- System.Void Hast::ExternalInvocationProxy() start
    \Finished\ <= \FinishedInternal\;
    \Hast::ExternalInvocationProxy()\: process (\Clock\) 
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \FinishedInternal\ <= false;
                \Hast::ExternalInvocationProxy().ParallelAlgorithm::Run(SimpleMemory)._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().ObjectOrientedShowcase::Run(SimpleMemory)._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumberAsync(SimpleMemory)._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().PrimeCalculator::ArePrimeNumbers(SimpleMemory)._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory)._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory)._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().RecursiveAlgorithms::CalculateFactorial(SimpleMemory)._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().SimdCalculator::AddVectors(SimpleMemory)._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().SimdCalculator::SubtractVectors(SimpleMemory)._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().SimdCalculator::MultiplyVectors(SimpleMemory)._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().SimdCalculator::DivideVectors(SimpleMemory)._Started.0\ <= false;
            else 
                if (\Started\ = true and \FinishedInternal\ = false) then 
                    -- Starting the state machine corresponding to the given member ID.
                    case \MemberId\ is 
                        when 0 => 
                            if (\Hast::ExternalInvocationProxy().ParallelAlgorithm::Run(SimpleMemory)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().ParallelAlgorithm::Run(SimpleMemory)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().ParallelAlgorithm::Run(SimpleMemory)._Started.0\ = \Hast::ExternalInvocationProxy().ParallelAlgorithm::Run(SimpleMemory)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().ParallelAlgorithm::Run(SimpleMemory)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 1 => 
                            if (\Hast::ExternalInvocationProxy().ObjectOrientedShowcase::Run(SimpleMemory)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().ObjectOrientedShowcase::Run(SimpleMemory)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().ObjectOrientedShowcase::Run(SimpleMemory)._Started.0\ = \Hast::ExternalInvocationProxy().ObjectOrientedShowcase::Run(SimpleMemory)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().ObjectOrientedShowcase::Run(SimpleMemory)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 2 => 
                            if (\Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\ = \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 3 => 
                            if (\Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumberAsync(SimpleMemory)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumberAsync(SimpleMemory)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumberAsync(SimpleMemory)._Started.0\ = \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumberAsync(SimpleMemory)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumberAsync(SimpleMemory)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 4 => 
                            if (\Hast::ExternalInvocationProxy().PrimeCalculator::ArePrimeNumbers(SimpleMemory)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().PrimeCalculator::ArePrimeNumbers(SimpleMemory)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().PrimeCalculator::ArePrimeNumbers(SimpleMemory)._Started.0\ = \Hast::ExternalInvocationProxy().PrimeCalculator::ArePrimeNumbers(SimpleMemory)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().PrimeCalculator::ArePrimeNumbers(SimpleMemory)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 5 => 
                            if (\Hast::ExternalInvocationProxy().PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory)._Started.0\ = \Hast::ExternalInvocationProxy().PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 6 => 
                            if (\Hast::ExternalInvocationProxy().RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory)._Started.0\ = \Hast::ExternalInvocationProxy().RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 7 => 
                            if (\Hast::ExternalInvocationProxy().RecursiveAlgorithms::CalculateFactorial(SimpleMemory)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().RecursiveAlgorithms::CalculateFactorial(SimpleMemory)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().RecursiveAlgorithms::CalculateFactorial(SimpleMemory)._Started.0\ = \Hast::ExternalInvocationProxy().RecursiveAlgorithms::CalculateFactorial(SimpleMemory)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().RecursiveAlgorithms::CalculateFactorial(SimpleMemory)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 8 => 
                            if (\Hast::ExternalInvocationProxy().SimdCalculator::AddVectors(SimpleMemory)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().SimdCalculator::AddVectors(SimpleMemory)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().SimdCalculator::AddVectors(SimpleMemory)._Started.0\ = \Hast::ExternalInvocationProxy().SimdCalculator::AddVectors(SimpleMemory)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().SimdCalculator::AddVectors(SimpleMemory)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 9 => 
                            if (\Hast::ExternalInvocationProxy().SimdCalculator::SubtractVectors(SimpleMemory)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().SimdCalculator::SubtractVectors(SimpleMemory)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().SimdCalculator::SubtractVectors(SimpleMemory)._Started.0\ = \Hast::ExternalInvocationProxy().SimdCalculator::SubtractVectors(SimpleMemory)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().SimdCalculator::SubtractVectors(SimpleMemory)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 10 => 
                            if (\Hast::ExternalInvocationProxy().SimdCalculator::MultiplyVectors(SimpleMemory)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().SimdCalculator::MultiplyVectors(SimpleMemory)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().SimdCalculator::MultiplyVectors(SimpleMemory)._Started.0\ = \Hast::ExternalInvocationProxy().SimdCalculator::MultiplyVectors(SimpleMemory)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().SimdCalculator::MultiplyVectors(SimpleMemory)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 11 => 
                            if (\Hast::ExternalInvocationProxy().SimdCalculator::DivideVectors(SimpleMemory)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().SimdCalculator::DivideVectors(SimpleMemory)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().SimdCalculator::DivideVectors(SimpleMemory)._Started.0\ = \Hast::ExternalInvocationProxy().SimdCalculator::DivideVectors(SimpleMemory)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().SimdCalculator::DivideVectors(SimpleMemory)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when others => 
                            null;
                    end case;
                else 
                    -- Waiting for Started to be pulled back to zero that signals the framework noting the finish.
                    if (\Started\ = false and \FinishedInternal\ = true) then 
                        \FinishedInternal\ <= false;
                    end if;
                end if;
            end if;
        end if;
    end process;
    -- System.Void Hast::ExternalInvocationProxy() end


    -- System.Void Hast::InternalInvocationProxy().System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32) start
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.ParallelAlgorithm::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 (#0):
    \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._Started\ <= \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.0\;
    \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.indexObject.parameter.In\ <= \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).indexObject.parameter.Out.0\;
    \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Finished.0\ <= \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0._Finished\;
    \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).return.0\ <= \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).0.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.ParallelAlgorithm::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 (#1):
    \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._Started\ <= \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.1\;
    \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.indexObject.parameter.In\ <= \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).indexObject.parameter.Out.1\;
    \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Finished.1\ <= \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1._Finished\;
    \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).return.1\ <= \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).1.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.ParallelAlgorithm::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 (#2):
    \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._Started\ <= \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.2\;
    \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.indexObject.parameter.In\ <= \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).indexObject.parameter.Out.2\;
    \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Finished.2\ <= \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2._Finished\;
    \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).return.2\ <= \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).2.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.ParallelAlgorithm::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 (#3):
    \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._Started\ <= \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.3\;
    \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.indexObject.parameter.In\ <= \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).indexObject.parameter.Out.3\;
    \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Finished.3\ <= \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3._Finished\;
    \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).return.3\ <= \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).3.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.ParallelAlgorithm::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 (#4):
    \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._Started\ <= \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Started.4\;
    \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.indexObject.parameter.In\ <= \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).indexObject.parameter.Out.4\;
    \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32)._Finished.4\ <= \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4._Finished\;
    \ParallelAlgorithm::Run(SimpleMemory).0.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).return.4\ <= \ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(UInt32).4.return\;
    -- System.Void Hast::InternalInvocationProxy().System.UInt32 Hast.Samples.SampleAssembly.ParallelAlgorithm/<>c__DisplayClass3_0::<Run>b__0(System.UInt32) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.MemoryContainer::.ctor(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) start
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.ObjectOrientedShowcase::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 (#0):
    \MemoryContainer::.ctor(SimpleMemory).0._Started\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::.ctor(SimpleMemory)._Started.0\;
    \MemoryContainer::.ctor(SimpleMemory).0.this.parameter.In\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::.ctor(SimpleMemory).this.parameter.Out.0\;
    \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::.ctor(SimpleMemory)._Finished.0\ <= \MemoryContainer::.ctor(SimpleMemory).0._Finished\;
    \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::.ctor(SimpleMemory).this.parameter.In.0\ <= \MemoryContainer::.ctor(SimpleMemory).0.this.parameter.Out\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.MemoryContainer::.ctor(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) end


    -- System.Void Hast::InternalInvocationProxy().System.UInt32 Hast.Samples.SampleAssembly.MemoryContainer::GetInput() start
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.ObjectOrientedShowcase::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 (#0):
    \MemoryContainer::GetInput().0._Started\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::GetInput()._Started.0\;
    \MemoryContainer::GetInput().0.this.parameter.In\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::GetInput().this.parameter.Out.0\;
    \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::GetInput()._Finished.0\ <= \MemoryContainer::GetInput().0._Finished\;
    \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::GetInput().return.0\ <= \MemoryContainer::GetInput().0.return\;
    \ObjectOrientedShowcase::Run(SimpleMemory).0.MemoryContainer::GetInput().this.parameter.In.0\ <= \MemoryContainer::GetInput().0.this.parameter.Out\;
    -- System.Void Hast::InternalInvocationProxy().System.UInt32 Hast.Samples.SampleAssembly.MemoryContainer::GetInput() end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.NumberContainer::.ctor() start
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.ObjectOrientedShowcase::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 (#0):
    \NumberContainer::.ctor().0._Started\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor()._Started.0\;
    \NumberContainer::.ctor().0.this.parameter.In\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor().this.parameter.Out.0\;
    \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor()._Finished.0\ <= \NumberContainer::.ctor().0._Finished\;
    \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor().this.parameter.In.0\ <= \NumberContainer::.ctor().0.this.parameter.Out\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.NumberContainer::.ctor() end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.NumberContainer::.ctor(System.UInt32) start
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.ObjectOrientedShowcase::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 (#0):
    \NumberContainer::.ctor(UInt32).0._Started\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor(UInt32)._Started.0\;
    \NumberContainer::.ctor(UInt32).0.this.parameter.In\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor(UInt32).this.parameter.Out.0\;
    \NumberContainer::.ctor(UInt32).0.number.parameter.In\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor(UInt32).number.parameter.Out.0\;
    \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor(UInt32)._Finished.0\ <= \NumberContainer::.ctor(UInt32).0._Finished\;
    \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::.ctor(UInt32).this.parameter.In.0\ <= \NumberContainer::.ctor(UInt32).0.this.parameter.Out\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.NumberContainer::.ctor(System.UInt32) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.NumberContainer::set_NumberPlusFive(System.UInt32) start
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.ObjectOrientedShowcase::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 (#0):
    \NumberContainer::set_NumberPlusFive(UInt32).0._Started\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::set_NumberPlusFive(UInt32)._Started.0\;
    \NumberContainer::set_NumberPlusFive(UInt32).0.this.parameter.In\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::set_NumberPlusFive(UInt32).this.parameter.Out.0\;
    \NumberContainer::set_NumberPlusFive(UInt32).0.value.parameter.In\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::set_NumberPlusFive(UInt32).value.parameter.Out.0\;
    \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::set_NumberPlusFive(UInt32)._Finished.0\ <= \NumberContainer::set_NumberPlusFive(UInt32).0._Finished\;
    \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::set_NumberPlusFive(UInt32).this.parameter.In.0\ <= \NumberContainer::set_NumberPlusFive(UInt32).0.this.parameter.Out\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.NumberContainer::set_NumberPlusFive(System.UInt32) end


    -- System.Void Hast::InternalInvocationProxy().System.UInt32 Hast.Samples.SampleAssembly.NumberContainer::IncreaseNumber(System.UInt32) start
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.ObjectOrientedShowcase::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 (#0):
    \NumberContainer::IncreaseNumber(UInt32).0._Started\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32)._Started.0\;
    \NumberContainer::IncreaseNumber(UInt32).0.this.parameter.In\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32).this.parameter.Out.0\;
    \NumberContainer::IncreaseNumber(UInt32).0.increaseBy.parameter.In\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32).increaseBy.parameter.Out.0\;
    \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32)._Finished.0\ <= \NumberContainer::IncreaseNumber(UInt32).0._Finished\;
    \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32).return.0\ <= \NumberContainer::IncreaseNumber(UInt32).0.return\;
    \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::IncreaseNumber(UInt32).this.parameter.In.0\ <= \NumberContainer::IncreaseNumber(UInt32).0.this.parameter.Out\;
    -- System.Void Hast::InternalInvocationProxy().System.UInt32 Hast.Samples.SampleAssembly.NumberContainer::IncreaseNumber(System.UInt32) end


    -- System.Void Hast::InternalInvocationProxy().System.UInt32 Hast.Samples.SampleAssembly.NumberContainer::get_NumberPlusFive() start
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.ObjectOrientedShowcase::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 (#0):
    \NumberContainer::get_NumberPlusFive().0._Started\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::get_NumberPlusFive()._Started.0\;
    \NumberContainer::get_NumberPlusFive().0.this.parameter.In\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::get_NumberPlusFive().this.parameter.Out.0\;
    \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::get_NumberPlusFive()._Finished.0\ <= \NumberContainer::get_NumberPlusFive().0._Finished\;
    \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::get_NumberPlusFive().return.0\ <= \NumberContainer::get_NumberPlusFive().0.return\;
    \ObjectOrientedShowcase::Run(SimpleMemory).0.NumberContainer::get_NumberPlusFive().this.parameter.In.0\ <= \NumberContainer::get_NumberPlusFive().0.this.parameter.Out\;
    -- System.Void Hast::InternalInvocationProxy().System.UInt32 Hast.Samples.SampleAssembly.NumberContainer::get_NumberPlusFive() end


    -- System.Void Hast::InternalInvocationProxy().System.UInt32 Hast.Samples.SampleAssembly.ObjectOrientedShowcase::SumNumberCointainers(Hast.Samples.SampleAssembly.NumberContainer[]) start
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.ObjectOrientedShowcase::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 (#0):
    \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._Started\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[])._Started.0\;
    \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.numberContainers.parameter.In\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).numberContainers.parameter.Out.0\;
    \ObjectOrientedShowcase::Run(SimpleMemory).0.ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[])._Finished.0\ <= \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0._Finished\;
    \ObjectOrientedShowcase::Run(SimpleMemory).0.ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).return.0\ <= \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.return\;
    \ObjectOrientedShowcase::Run(SimpleMemory).0.ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).numberContainers.parameter.In.0\ <= \ObjectOrientedShowcase::SumNumberCointainers(NumberContainer[]).0.numberContainers.parameter.Out\;
    -- System.Void Hast::InternalInvocationProxy().System.UInt32 Hast.Samples.SampleAssembly.ObjectOrientedShowcase::SumNumberCointainers(Hast.Samples.SampleAssembly.NumberContainer[]) end


    -- System.Void Hast::InternalInvocationProxy().System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberInternal(System.UInt32) start
    \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\ <= false;
                \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.Void Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumber(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0
                case \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\) then 
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.runningIndex.0\ := 0;
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Started\ <= true;
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.number.parameter.In\ <= \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).number.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.runningIndex.0\ is 
                            when 0 => 
                                if (\PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\ <= true;
                                    \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Started\ <= false;
                                    \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).return.0\ <= \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::IsPrimeNumber(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ArePrimeNumbers(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0
                case \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\) then 
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.runningIndex.0\ := 0;
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Started\ <= true;
                            \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.number.parameter.In\ <= \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).number.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.runningIndex.0\ is 
                            when 0 => 
                                if (\PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\ <= true;
                                    \PrimeCalculator::IsPrimeNumberInternal(UInt32).0._Started\ <= false;
                                    \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32).return.0\ <= \PrimeCalculator::IsPrimeNumberInternal(UInt32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumberInternal(UInt32).PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                            \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.PrimeCalculator::IsPrimeNumberInternal(UInt32)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberInternal(System.UInt32) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumber(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) start
    \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).Hast::ExternalInvocationProxy().runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).Hast::ExternalInvocationProxy().runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).Hast::ExternalInvocationProxy().runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).Hast::ExternalInvocationProxy().runningState.0\ := WaitingForStarted;
                \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\ <= false;
                \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.Threading.Tasks.Task Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberAsync(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0
                case \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\) then 
                            \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.runningIndex.0\ := 0;
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Started\ <= true;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.runningIndex.0\ is 
                            when 0 => 
                                if (\PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\ <= true;
                                    \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Started\ <= false;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                            \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0.PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Void Hast::ExternalInvocationProxy()
                case \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).Hast::ExternalInvocationProxy().runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\) then 
                            \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).Hast::ExternalInvocationProxy().runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).Hast::ExternalInvocationProxy().runningIndex.0\ := 0;
                            \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Started\ <= true;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).Hast::ExternalInvocationProxy().runningIndex.0\ is 
                            when 0 => 
                                if (\PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).Hast::ExternalInvocationProxy().runningState.0\ := AfterFinished;
                                    \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\ <= true;
                                    \PrimeCalculator::IsPrimeNumber(SimpleMemory).0._Started\ <= false;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory).Hast::ExternalInvocationProxy().runningState.0\ := WaitingForStarted;
                            \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumber(SimpleMemory)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumber(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) end


    -- System.Void Hast::InternalInvocationProxy().System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32) start
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 (#0):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.0\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.numberObject.parameter.In\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).numberObject.parameter.Out.0\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Finished.0\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).return.0\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).0.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 (#1):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.1\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.numberObject.parameter.In\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).numberObject.parameter.Out.1\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Finished.1\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).return.1\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).1.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 (#2):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.2\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.numberObject.parameter.In\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).numberObject.parameter.Out.2\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Finished.2\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).return.2\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).2.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 (#3):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.3\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.numberObject.parameter.In\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).numberObject.parameter.Out.3\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Finished.3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).return.3\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).3.return\;
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 (#4):
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._Started\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Started.4\;
    \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.numberObject.parameter.In\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).numberObject.parameter.Out.4\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32)._Finished.4\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4._Finished\;
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).return.4\ <= \PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(UInt32).4.return\;
    -- System.Void Hast::InternalInvocationProxy().System.Boolean Hast.Samples.SampleAssembly.PrimeCalculator/<>c::<ParallelizedArePrimeNumbers>b__9_0(System.UInt32) end


    -- System.Void Hast::InternalInvocationProxy().System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16) start
    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\: \InternalInvocationProxy_boolean_Array\(5 downto 0) := (others => false);
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningIndex.0\: integer range 0 to 5 := 0;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.runningIndex.0\: integer range 0 to 5 := 0;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.runningIndex.0\: integer range 0 to 5 := 0;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.runningIndex.0\: integer range 0 to 5 := 0;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.runningIndex.0\: integer range 0 to 5 := 0;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.runningIndex.0\: integer range 0 to 5 := 0;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.runningIndex.0\: integer range 0 to 5 := 0;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\ := (others => false);
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.runningState.0\ := WaitingForStarted;
                \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= false;
            else 
                -- Building a boolean array where each of the elements will indicate whether the component with the given index should be started next.
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(0) := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Started\ = false;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(1) := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Started\ = false;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(2) := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Started\ = false;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(3) := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Started\ = false;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(4) := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Started\ = false;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(5) := \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Started\ = false;

                -- Invocation handler #0 out of 1 corresponding to System.Void Hast.Samples.SampleAssembly.RecursiveAlgorithms::CalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0
                case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\) then 
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= false;
                            case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\ is 
                                when (false, false, false, false, false, true) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningIndex.0\ := 0;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(0) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.number.parameter.In\ <= \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, false, true, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningIndex.0\ := 1;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(1) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.number.parameter.In\ <= \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, true, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningIndex.0\ := 2;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(2) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.number.parameter.In\ <= \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, true, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningIndex.0\ := 3;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(3) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.number.parameter.In\ <= \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, true, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningIndex.0\ := 4;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(4) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.number.parameter.In\ <= \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (true, false, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningIndex.0\ := 5;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(5) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.number.parameter.In\ <= \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when others => 
                                    null;
                            end case;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningIndex.0\ is 
                            when 0 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Started\ <= false;
                                    \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.return\;
                                end if;
                            when 1 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Started\ <= false;
                                    \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.return\;
                                end if;
                            when 2 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Started\ <= false;
                                    \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.return\;
                                end if;
                            when 3 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Started\ <= false;
                                    \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.return\;
                                end if;
                            when 4 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Started\ <= false;
                                    \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.return\;
                                end if;
                            when 5 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Started\ <= false;
                                    \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                            \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).0
                case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= false;
                            case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\ is 
                                when (false, false, false, false, false, true) => 
                                    -- The component can't invoke itself, so not putting anything here.
                                    null;
                                when (false, false, false, false, true, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.runningIndex.0\ := 1;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(1) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, true, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.runningIndex.0\ := 2;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(2) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, true, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.runningIndex.0\ := 3;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(3) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, true, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.runningIndex.0\ := 4;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(4) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (true, false, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.runningIndex.0\ := 5;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(5) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when others => 
                                    null;
                            end case;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.runningIndex.0\ is 
                            when 0 => 
                                -- The component can't invoke itself, so not putting anything here.
                                null;
                            when 1 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.return\;
                                end if;
                            when 2 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.return\;
                                end if;
                            when 3 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.return\;
                                end if;
                            when 4 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.return\;
                                end if;
                            when 5 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.runningState.0\ := WaitingForStarted;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).1
                case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= false;
                            case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\ is 
                                when (false, false, false, false, false, true) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.runningIndex.0\ := 0;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(0) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, false, true, false) => 
                                    -- The component can't invoke itself, so not putting anything here.
                                    null;
                                when (false, false, false, true, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.runningIndex.0\ := 2;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(2) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, true, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.runningIndex.0\ := 3;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(3) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, true, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.runningIndex.0\ := 4;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(4) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (true, false, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.runningIndex.0\ := 5;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(5) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when others => 
                                    null;
                            end case;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.runningIndex.0\ is 
                            when 0 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.return\;
                                end if;
                            when 1 => 
                                -- The component can't invoke itself, so not putting anything here.
                                null;
                            when 2 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.return\;
                                end if;
                            when 3 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.return\;
                                end if;
                            when 4 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.return\;
                                end if;
                            when 5 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.runningState.0\ := WaitingForStarted;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).2
                case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= false;
                            case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\ is 
                                when (false, false, false, false, false, true) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.runningIndex.0\ := 0;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(0) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, false, true, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.runningIndex.0\ := 1;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(1) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, true, false, false) => 
                                    -- The component can't invoke itself, so not putting anything here.
                                    null;
                                when (false, false, true, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.runningIndex.0\ := 3;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(3) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, true, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.runningIndex.0\ := 4;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(4) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (true, false, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.runningIndex.0\ := 5;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(5) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when others => 
                                    null;
                            end case;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.runningIndex.0\ is 
                            when 0 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.return\;
                                end if;
                            when 1 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.return\;
                                end if;
                            when 2 => 
                                -- The component can't invoke itself, so not putting anything here.
                                null;
                            when 3 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.return\;
                                end if;
                            when 4 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.return\;
                                end if;
                            when 5 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.runningState.0\ := WaitingForStarted;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).3
                case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= false;
                            case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\ is 
                                when (false, false, false, false, false, true) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.runningIndex.0\ := 0;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(0) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, false, true, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.runningIndex.0\ := 1;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(1) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, true, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.runningIndex.0\ := 2;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(2) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, true, false, false, false) => 
                                    -- The component can't invoke itself, so not putting anything here.
                                    null;
                                when (false, true, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.runningIndex.0\ := 4;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(4) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (true, false, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.runningIndex.0\ := 5;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(5) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when others => 
                                    null;
                            end case;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.runningIndex.0\ is 
                            when 0 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.return\;
                                end if;
                            when 1 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.return\;
                                end if;
                            when 2 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.return\;
                                end if;
                            when 3 => 
                                -- The component can't invoke itself, so not putting anything here.
                                null;
                            when 4 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.return\;
                                end if;
                            when 5 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.runningState.0\ := WaitingForStarted;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).4
                case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= false;
                            case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\ is 
                                when (false, false, false, false, false, true) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.runningIndex.0\ := 0;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(0) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, false, true, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.runningIndex.0\ := 1;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(1) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, true, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.runningIndex.0\ := 2;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(2) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, true, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.runningIndex.0\ := 3;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(3) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, true, false, false, false, false) => 
                                    -- The component can't invoke itself, so not putting anything here.
                                    null;
                                when (true, false, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.runningIndex.0\ := 5;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(5) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when others => 
                                    null;
                            end case;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.runningIndex.0\ is 
                            when 0 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.return\;
                                end if;
                            when 1 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.return\;
                                end if;
                            when 2 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.return\;
                                end if;
                            when 3 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.return\;
                                end if;
                            when 4 => 
                                -- The component can't invoke itself, so not putting anything here.
                                null;
                            when 5 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.runningState.0\ := WaitingForStarted;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).5
                case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= false;
                            case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\ is 
                                when (false, false, false, false, false, true) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.runningIndex.0\ := 0;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(0) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, false, true, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.runningIndex.0\ := 1;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(1) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, true, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.runningIndex.0\ := 2;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(2) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, true, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.runningIndex.0\ := 3;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(3) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, true, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.runningIndex.0\ := 4;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).targetAvailableIndicator\(4) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (true, false, false, false, false, false) => 
                                    -- The component can't invoke itself, so not putting anything here.
                                    null;
                                when others => 
                                    null;
                            end case;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.runningIndex.0\ is 
                            when 0 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.return\;
                                end if;
                            when 1 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.return\;
                                end if;
                            when 2 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.return\;
                                end if;
                            when 3 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.return\;
                                end if;
                            when 4 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.return\;
                                end if;
                            when 5 => 
                                -- The component can't invoke itself, so not putting anything here.
                                null;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.runningState.0\ := WaitingForStarted;
                            \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16) end


    -- System.Void Hast::InternalInvocationProxy().System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16) start
    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\: \InternalInvocationProxy_boolean_Array\(5 downto 0) := (others => false);
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningIndex.0\: integer range 0 to 5 := 0;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.runningIndex.0\: integer range 0 to 5 := 0;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.runningIndex.0\: integer range 0 to 5 := 0;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.runningIndex.0\: integer range 0 to 5 := 0;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.runningIndex.0\: integer range 0 to 5 := 0;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.runningIndex.0\: integer range 0 to 5 := 0;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.runningIndex.0\: integer range 0 to 5 := 0;
        Variable \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\ := (others => false);
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.runningState.0\ := WaitingForStarted;
                \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= false;
                \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= false;
            else 
                -- Building a boolean array where each of the elements will indicate whether the component with the given index should be started next.
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(0) := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Started\ = false;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(1) := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Started\ = false;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(2) := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Started\ = false;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(3) := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Started\ = false;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(4) := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Started\ = true and \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Started\ = false;
                \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(5) := \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Started\ = false;

                -- Invocation handler #0 out of 1 corresponding to System.Void Hast.Samples.SampleAssembly.RecursiveAlgorithms::CalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0
                case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\) then 
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= false;
                            case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\ is 
                                when (false, false, false, false, false, true) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningIndex.0\ := 0;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(0) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.number.parameter.In\ <= \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, false, true, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningIndex.0\ := 1;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(1) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.number.parameter.In\ <= \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, true, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningIndex.0\ := 2;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(2) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.number.parameter.In\ <= \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, true, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningIndex.0\ := 3;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(3) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.number.parameter.In\ <= \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, true, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningIndex.0\ := 4;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(4) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.number.parameter.In\ <= \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (true, false, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningIndex.0\ := 5;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(5) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.number.parameter.In\ <= \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when others => 
                                    null;
                            end case;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningIndex.0\ is 
                            when 0 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Started\ <= false;
                                    \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.return\;
                                end if;
                            when 1 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Started\ <= false;
                                    \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.return\;
                                end if;
                            when 2 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Started\ <= false;
                                    \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.return\;
                                end if;
                            when 3 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Started\ <= false;
                                    \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.return\;
                                end if;
                            when 4 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Started\ <= false;
                                    \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.return\;
                                end if;
                            when 5 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Started\ <= false;
                                    \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                            \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).0
                case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= false;
                            case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\ is 
                                when (false, false, false, false, false, true) => 
                                    -- The component can't invoke itself, so not putting anything here.
                                    null;
                                when (false, false, false, false, true, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.runningIndex.0\ := 1;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(1) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, true, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.runningIndex.0\ := 2;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(2) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, true, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.runningIndex.0\ := 3;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(3) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, true, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.runningIndex.0\ := 4;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(4) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (true, false, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.runningIndex.0\ := 5;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(5) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when others => 
                                    null;
                            end case;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.runningIndex.0\ is 
                            when 0 => 
                                -- The component can't invoke itself, so not putting anything here.
                                null;
                            when 1 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.return\;
                                end if;
                            when 2 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.return\;
                                end if;
                            when 3 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.return\;
                                end if;
                            when 4 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.return\;
                                end if;
                            when 5 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.runningState.0\ := WaitingForStarted;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).1
                case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= false;
                            case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\ is 
                                when (false, false, false, false, false, true) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.runningIndex.0\ := 0;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(0) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, false, true, false) => 
                                    -- The component can't invoke itself, so not putting anything here.
                                    null;
                                when (false, false, false, true, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.runningIndex.0\ := 2;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(2) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, true, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.runningIndex.0\ := 3;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(3) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, true, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.runningIndex.0\ := 4;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(4) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (true, false, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.runningIndex.0\ := 5;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(5) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when others => 
                                    null;
                            end case;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.runningIndex.0\ is 
                            when 0 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.return\;
                                end if;
                            when 1 => 
                                -- The component can't invoke itself, so not putting anything here.
                                null;
                            when 2 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.return\;
                                end if;
                            when 3 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.return\;
                                end if;
                            when 4 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.return\;
                                end if;
                            when 5 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.runningState.0\ := WaitingForStarted;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).2
                case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= false;
                            case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\ is 
                                when (false, false, false, false, false, true) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.runningIndex.0\ := 0;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(0) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, false, true, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.runningIndex.0\ := 1;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(1) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, true, false, false) => 
                                    -- The component can't invoke itself, so not putting anything here.
                                    null;
                                when (false, false, true, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.runningIndex.0\ := 3;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(3) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, true, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.runningIndex.0\ := 4;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(4) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (true, false, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.runningIndex.0\ := 5;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(5) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when others => 
                                    null;
                            end case;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.runningIndex.0\ is 
                            when 0 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.return\;
                                end if;
                            when 1 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.return\;
                                end if;
                            when 2 => 
                                -- The component can't invoke itself, so not putting anything here.
                                null;
                            when 3 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.return\;
                                end if;
                            when 4 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.return\;
                                end if;
                            when 5 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.runningState.0\ := WaitingForStarted;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).3
                case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= false;
                            case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\ is 
                                when (false, false, false, false, false, true) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.runningIndex.0\ := 0;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(0) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, false, true, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.runningIndex.0\ := 1;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(1) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, true, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.runningIndex.0\ := 2;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(2) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, true, false, false, false) => 
                                    -- The component can't invoke itself, so not putting anything here.
                                    null;
                                when (false, true, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.runningIndex.0\ := 4;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(4) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (true, false, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.runningIndex.0\ := 5;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(5) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when others => 
                                    null;
                            end case;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.runningIndex.0\ is 
                            when 0 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.return\;
                                end if;
                            when 1 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.return\;
                                end if;
                            when 2 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.return\;
                                end if;
                            when 3 => 
                                -- The component can't invoke itself, so not putting anything here.
                                null;
                            when 4 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.return\;
                                end if;
                            when 5 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.runningState.0\ := WaitingForStarted;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).4
                case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= false;
                            case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\ is 
                                when (false, false, false, false, false, true) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.runningIndex.0\ := 0;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(0) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, false, true, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.runningIndex.0\ := 1;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(1) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, true, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.runningIndex.0\ := 2;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(2) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, true, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.runningIndex.0\ := 3;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(3) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, true, false, false, false, false) => 
                                    -- The component can't invoke itself, so not putting anything here.
                                    null;
                                when (true, false, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.runningIndex.0\ := 5;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(5) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when others => 
                                    null;
                            end case;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.runningIndex.0\ is 
                            when 0 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.return\;
                                end if;
                            when 1 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.return\;
                                end if;
                            when 2 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.return\;
                                end if;
                            when 3 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.return\;
                                end if;
                            when 4 => 
                                -- The component can't invoke itself, so not putting anything here.
                                null;
                            when 5 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.runningState.0\ := WaitingForStarted;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16).5
                case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\) then 
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= false;
                            case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\ is 
                                when (false, false, false, false, false, true) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.runningIndex.0\ := 0;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(0) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, false, true, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.runningIndex.0\ := 1;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(1) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, false, true, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.runningIndex.0\ := 2;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(2) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, false, true, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.runningIndex.0\ := 3;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(3) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (false, true, false, false, false, false) => 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.runningState.0\ := WaitingForFinished;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.runningIndex.0\ := 4;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Started\ <= true;
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).targetAvailableIndicator\(4) := false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.number.parameter.In\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).number.parameter.Out.0\;
                                when (true, false, false, false, false, false) => 
                                    -- The component can't invoke itself, so not putting anything here.
                                    null;
                                when others => 
                                    null;
                            end case;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.runningIndex.0\ is 
                            when 0 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.return\;
                                end if;
                            when 1 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.return\;
                                end if;
                            when 2 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.return\;
                                end if;
                            when 3 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.return\;
                                end if;
                            when 4 => 
                                if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Finished\) then 
                                    \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.runningState.0\ := AfterFinished;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= true;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4._Started\ <= false;
                                    \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).return.0\ <= \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.return\;
                                end if;
                            when 5 => 
                                -- The component can't invoke itself, so not putting anything here.
                                null;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.runningState.0\ := WaitingForStarted;
                            \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.UInt32 Hast.Samples.SampleAssembly.RecursiveAlgorithms::RecursivelyCalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,System.Int16) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.SimdCalculator::RunSimdOperation(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,Hast.Samples.SampleAssembly.SimdOperation) start
    \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::AddVectors(SimpleMemory).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::AddVectors(SimpleMemory).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::SubtractVectors(SimpleMemory).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::SubtractVectors(SimpleMemory).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::MultiplyVectors(SimpleMemory).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::MultiplyVectors(SimpleMemory).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::DivideVectors(SimpleMemory).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::DivideVectors(SimpleMemory).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::AddVectors(SimpleMemory).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::AddVectors(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::SubtractVectors(SimpleMemory).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::SubtractVectors(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::MultiplyVectors(SimpleMemory).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::MultiplyVectors(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::DivideVectors(SimpleMemory).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::DivideVectors(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                \SimdCalculator::AddVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\ <= false;
                \SimdCalculator::SubtractVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\ <= false;
                \SimdCalculator::MultiplyVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\ <= false;
                \SimdCalculator::DivideVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.Void Hast.Samples.SampleAssembly.SimdCalculator::AddVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0
                case \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::AddVectors(SimpleMemory).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\SimdCalculator::AddVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\) then 
                            \SimdCalculator::AddVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::AddVectors(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::AddVectors(SimpleMemory).0.runningIndex.0\ := 0;
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._Started\ <= true;
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.operation.parameter.In\ <= \SimdCalculator::AddVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).operation.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::AddVectors(SimpleMemory).0.runningIndex.0\ is 
                            when 0 => 
                                if (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::AddVectors(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \SimdCalculator::AddVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\ <= true;
                                    \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._Started\ <= false;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\SimdCalculator::AddVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::AddVectors(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                            \SimdCalculator::AddVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Void Hast.Samples.SampleAssembly.SimdCalculator::SubtractVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0
                case \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::SubtractVectors(SimpleMemory).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\SimdCalculator::SubtractVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\) then 
                            \SimdCalculator::SubtractVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::SubtractVectors(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::SubtractVectors(SimpleMemory).0.runningIndex.0\ := 0;
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._Started\ <= true;
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.operation.parameter.In\ <= \SimdCalculator::SubtractVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).operation.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::SubtractVectors(SimpleMemory).0.runningIndex.0\ is 
                            when 0 => 
                                if (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::SubtractVectors(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \SimdCalculator::SubtractVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\ <= true;
                                    \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._Started\ <= false;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\SimdCalculator::SubtractVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::SubtractVectors(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                            \SimdCalculator::SubtractVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Void Hast.Samples.SampleAssembly.SimdCalculator::MultiplyVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0
                case \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::MultiplyVectors(SimpleMemory).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\SimdCalculator::MultiplyVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\) then 
                            \SimdCalculator::MultiplyVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::MultiplyVectors(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::MultiplyVectors(SimpleMemory).0.runningIndex.0\ := 0;
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._Started\ <= true;
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.operation.parameter.In\ <= \SimdCalculator::MultiplyVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).operation.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::MultiplyVectors(SimpleMemory).0.runningIndex.0\ is 
                            when 0 => 
                                if (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::MultiplyVectors(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \SimdCalculator::MultiplyVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\ <= true;
                                    \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._Started\ <= false;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\SimdCalculator::MultiplyVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::MultiplyVectors(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                            \SimdCalculator::MultiplyVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Void Hast.Samples.SampleAssembly.SimdCalculator::DivideVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0
                case \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::DivideVectors(SimpleMemory).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\SimdCalculator::DivideVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\) then 
                            \SimdCalculator::DivideVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::DivideVectors(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::DivideVectors(SimpleMemory).0.runningIndex.0\ := 0;
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._Started\ <= true;
                            \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.operation.parameter.In\ <= \SimdCalculator::DivideVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).operation.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::DivideVectors(SimpleMemory).0.runningIndex.0\ is 
                            when 0 => 
                                if (\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::DivideVectors(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \SimdCalculator::DivideVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\ <= true;
                                    \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0._Started\ <= false;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\SimdCalculator::DivideVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).SimdCalculator::DivideVectors(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                            \SimdCalculator::DivideVectors(SimpleMemory).0.SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.SimdCalculator::RunSimdOperation(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory,Hast.Samples.SampleAssembly.SimdOperation) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.ParallelAlgorithm::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \ParallelAlgorithm::Run(SimpleMemory).0._Started\ <= \Hast::ExternalInvocationProxy().ParallelAlgorithm::Run(SimpleMemory)._Started.0\;
    \Hast::ExternalInvocationProxy().ParallelAlgorithm::Run(SimpleMemory)._Finished.0\ <= \ParallelAlgorithm::Run(SimpleMemory).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.ParallelAlgorithm::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.ObjectOrientedShowcase::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \ObjectOrientedShowcase::Run(SimpleMemory).0._Started\ <= \Hast::ExternalInvocationProxy().ObjectOrientedShowcase::Run(SimpleMemory)._Started.0\;
    \Hast::ExternalInvocationProxy().ObjectOrientedShowcase::Run(SimpleMemory)._Finished.0\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.ObjectOrientedShowcase::Run(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) end


    -- System.Void Hast::InternalInvocationProxy().System.Threading.Tasks.Task Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberAsync(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._Started\ <= \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumberAsync(SimpleMemory)._Started.0\;
    \Hast::ExternalInvocationProxy().PrimeCalculator::IsPrimeNumberAsync(SimpleMemory)._Finished.0\ <= \PrimeCalculator::IsPrimeNumberAsync(SimpleMemory).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Threading.Tasks.Task Hast.Samples.SampleAssembly.PrimeCalculator::IsPrimeNumberAsync(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ArePrimeNumbers(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._Started\ <= \Hast::ExternalInvocationProxy().PrimeCalculator::ArePrimeNumbers(SimpleMemory)._Started.0\;
    \Hast::ExternalInvocationProxy().PrimeCalculator::ArePrimeNumbers(SimpleMemory)._Finished.0\ <= \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ArePrimeNumbers(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._Started\ <= \Hast::ExternalInvocationProxy().PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory)._Started.0\;
    \Hast::ExternalInvocationProxy().PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory)._Finished.0\ <= \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.PrimeCalculator::ParallelizedArePrimeNumbers(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.RecursiveAlgorithms::CalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._Started\ <= \Hast::ExternalInvocationProxy().RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory)._Started.0\;
    \Hast::ExternalInvocationProxy().RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory)._Finished.0\ <= \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.RecursiveAlgorithms::CalculateFibonacchiSeries(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.RecursiveAlgorithms::CalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._Started\ <= \Hast::ExternalInvocationProxy().RecursiveAlgorithms::CalculateFactorial(SimpleMemory)._Started.0\;
    \Hast::ExternalInvocationProxy().RecursiveAlgorithms::CalculateFactorial(SimpleMemory)._Finished.0\ <= \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.RecursiveAlgorithms::CalculateFactorial(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.SimdCalculator::AddVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \SimdCalculator::AddVectors(SimpleMemory).0._Started\ <= \Hast::ExternalInvocationProxy().SimdCalculator::AddVectors(SimpleMemory)._Started.0\;
    \Hast::ExternalInvocationProxy().SimdCalculator::AddVectors(SimpleMemory)._Finished.0\ <= \SimdCalculator::AddVectors(SimpleMemory).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.SimdCalculator::AddVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.SimdCalculator::SubtractVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \SimdCalculator::SubtractVectors(SimpleMemory).0._Started\ <= \Hast::ExternalInvocationProxy().SimdCalculator::SubtractVectors(SimpleMemory)._Started.0\;
    \Hast::ExternalInvocationProxy().SimdCalculator::SubtractVectors(SimpleMemory)._Finished.0\ <= \SimdCalculator::SubtractVectors(SimpleMemory).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.SimdCalculator::SubtractVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.SimdCalculator::MultiplyVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \SimdCalculator::MultiplyVectors(SimpleMemory).0._Started\ <= \Hast::ExternalInvocationProxy().SimdCalculator::MultiplyVectors(SimpleMemory)._Started.0\;
    \Hast::ExternalInvocationProxy().SimdCalculator::MultiplyVectors(SimpleMemory)._Finished.0\ <= \SimdCalculator::MultiplyVectors(SimpleMemory).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.SimdCalculator::MultiplyVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.SimdCalculator::DivideVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \SimdCalculator::DivideVectors(SimpleMemory).0._Started\ <= \Hast::ExternalInvocationProxy().SimdCalculator::DivideVectors(SimpleMemory)._Started.0\;
    \Hast::ExternalInvocationProxy().SimdCalculator::DivideVectors(SimpleMemory)._Finished.0\ <= \SimdCalculator::DivideVectors(SimpleMemory).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.SimdCalculator::DivideVectors(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) end


    -- System.Void Hast::SimpleMemoryOperationProxy() start
    \CellIndex\ <= to_integer(\ParallelAlgorithm::Run(SimpleMemory).0.SimpleMemory.CellIndex\) when \ParallelAlgorithm::Run(SimpleMemory).0.SimpleMemory.ReadEnable\ or \ParallelAlgorithm::Run(SimpleMemory).0.SimpleMemory.WriteEnable\ else to_integer(\ObjectOrientedShowcase::Run(SimpleMemory).0.SimpleMemory.CellIndex\) when \ObjectOrientedShowcase::Run(SimpleMemory).0.SimpleMemory.ReadEnable\ or \ObjectOrientedShowcase::Run(SimpleMemory).0.SimpleMemory.WriteEnable\ else to_integer(\MemoryContainer::GetInput().0.SimpleMemory.CellIndex\) when \MemoryContainer::GetInput().0.SimpleMemory.ReadEnable\ or \MemoryContainer::GetInput().0.SimpleMemory.WriteEnable\ else to_integer(\PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.CellIndex\) when \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.ReadEnable\ or \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.WriteEnable\ else to_integer(\PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.CellIndex\) when \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ or \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ else to_integer(\PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.CellIndex\) when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ or \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ else to_integer(\RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.CellIndex\) when \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.WriteEnable\ else to_integer(\RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.CellIndex\) when \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.WriteEnable\ else to_integer(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.SimpleMemory.CellIndex\) when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.SimpleMemory.WriteEnable\ else to_integer(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.SimpleMemory.CellIndex\) when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.SimpleMemory.WriteEnable\ else to_integer(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.SimpleMemory.CellIndex\) when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.SimpleMemory.WriteEnable\ else to_integer(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.SimpleMemory.CellIndex\) when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.SimpleMemory.WriteEnable\ else to_integer(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.SimpleMemory.CellIndex\) when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.SimpleMemory.WriteEnable\ else to_integer(\RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.SimpleMemory.CellIndex\) when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.SimpleMemory.WriteEnable\ else to_integer(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.SimpleMemory.CellIndex\) when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.SimpleMemory.WriteEnable\ else to_integer(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.SimpleMemory.CellIndex\) when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.SimpleMemory.WriteEnable\ else to_integer(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.SimpleMemory.CellIndex\) when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.SimpleMemory.WriteEnable\ else to_integer(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.SimpleMemory.CellIndex\) when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.SimpleMemory.WriteEnable\ else to_integer(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.SimpleMemory.CellIndex\) when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.SimpleMemory.WriteEnable\ else to_integer(\RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.SimpleMemory.CellIndex\) when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.SimpleMemory.WriteEnable\ else to_integer(\SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.CellIndex\) when \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.ReadEnable\ or \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.WriteEnable\ else 0;
    \DataOut\ <= \ParallelAlgorithm::Run(SimpleMemory).0.SimpleMemory.DataOut\ when \ParallelAlgorithm::Run(SimpleMemory).0.SimpleMemory.WriteEnable\ else \ObjectOrientedShowcase::Run(SimpleMemory).0.SimpleMemory.DataOut\ when \ObjectOrientedShowcase::Run(SimpleMemory).0.SimpleMemory.WriteEnable\ else \MemoryContainer::GetInput().0.SimpleMemory.DataOut\ when \MemoryContainer::GetInput().0.SimpleMemory.WriteEnable\ else \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.DataOut\ when \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.WriteEnable\ else \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.DataOut\ when \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ else \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.DataOut\ when \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ else \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.DataOut\ when \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.WriteEnable\ else \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.DataOut\ when \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.WriteEnable\ else \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.SimpleMemory.DataOut\ when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.SimpleMemory.WriteEnable\ else \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.SimpleMemory.DataOut\ when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.SimpleMemory.WriteEnable\ else \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.SimpleMemory.DataOut\ when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.SimpleMemory.WriteEnable\ else \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.SimpleMemory.DataOut\ when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.SimpleMemory.WriteEnable\ else \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.SimpleMemory.DataOut\ when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.SimpleMemory.WriteEnable\ else \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.SimpleMemory.DataOut\ when \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.SimpleMemory.WriteEnable\ else \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.SimpleMemory.DataOut\ when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.SimpleMemory.WriteEnable\ else \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.SimpleMemory.DataOut\ when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.SimpleMemory.WriteEnable\ else \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.SimpleMemory.DataOut\ when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.SimpleMemory.WriteEnable\ else \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.SimpleMemory.DataOut\ when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.SimpleMemory.WriteEnable\ else \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.SimpleMemory.DataOut\ when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.SimpleMemory.WriteEnable\ else \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.SimpleMemory.DataOut\ when \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.SimpleMemory.WriteEnable\ else \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.DataOut\ when \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.WriteEnable\ else "00000000000000000000000000000000";
    \ReadEnable\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.SimpleMemory.ReadEnable\ or \MemoryContainer::GetInput().0.SimpleMemory.ReadEnable\ or \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.ReadEnable\ or \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ or \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.SimpleMemory.ReadEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.SimpleMemory.ReadEnable\ or \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.ReadEnable\ or \ParallelAlgorithm::Run(SimpleMemory).0.SimpleMemory.ReadEnable\;
    \WriteEnable\ <= \ObjectOrientedShowcase::Run(SimpleMemory).0.SimpleMemory.WriteEnable\ or \MemoryContainer::GetInput().0.SimpleMemory.WriteEnable\ or \PrimeCalculator::IsPrimeNumber(SimpleMemory).0.SimpleMemory.WriteEnable\ or \PrimeCalculator::ArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ or \PrimeCalculator::ParallelizedArePrimeNumbers(SimpleMemory).0.SimpleMemory.WriteEnable\ or \RecursiveAlgorithms::CalculateFibonacchiSeries(SimpleMemory).0.SimpleMemory.WriteEnable\ or \RecursiveAlgorithms::CalculateFactorial(SimpleMemory).0.SimpleMemory.WriteEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).0.SimpleMemory.WriteEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).1.SimpleMemory.WriteEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).2.SimpleMemory.WriteEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).3.SimpleMemory.WriteEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).4.SimpleMemory.WriteEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFibonacchiSeries(SimpleMemory,Int16).5.SimpleMemory.WriteEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).0.SimpleMemory.WriteEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).1.SimpleMemory.WriteEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).2.SimpleMemory.WriteEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).3.SimpleMemory.WriteEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).4.SimpleMemory.WriteEnable\ or \RecursiveAlgorithms::RecursivelyCalculateFactorial(SimpleMemory,Int16).5.SimpleMemory.WriteEnable\ or \SimdCalculator::RunSimdOperation(SimpleMemory,SimdOperation).0.SimpleMemory.WriteEnable\ or \ParallelAlgorithm::Run(SimpleMemory).0.SimpleMemory.WriteEnable\;
    -- System.Void Hast::SimpleMemoryOperationProxy() end

end Imp;
