library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library Hast;
use Hast.SimpleMemory.all;

entity Hast_IP is 
    port(
        \DataIn\: In std_logic_vector(31 downto 0);
        \DataOut\: Out std_logic_vector(31 downto 0);
        \CellIndex\: Out integer;
        \ReadEnable\: Out boolean;
        \WriteEnable\: Out boolean;
        \ReadsDone\: In boolean;
        \WritesDone\: In boolean;
        \MemberId\: In integer;
        \Reset\: In std_logic;
        \Started\: In boolean;
        \Finished\: Out boolean;
        \Clock\: In std_logic
    );
    -- Hast_IP ID: e1bfe8bd0d5d2e19934a8b929e75f51c7421cc348a2a84fd92bc0ad4cba032ac
    -- (Date and time removed for approval testing.)
    -- Generated by Hastlayer - hastlayer.com
end Hast_IP;

architecture Imp of Hast_IP is 
    -- This IP was generated by Hastlayer from .NET code to mimic the original logic. Note the following:
    -- * For each member (methods, functions) in .NET a state machine was generated. Each state machine's name corresponds to 
    --   the original member's name.
    -- * Inputs and outputs are passed between state machines as shared objects.
    -- * There are operations that take multiple clock cycles like interacting with the memory and long-running arithmetic operations 
    --   (modulo, division, multiplication). These are awaited in subsequent states but be aware that some states can take more 
    --   than one clock cycle to produce their output.
    -- * The ExternalInvocationProxy process dispatches invocations that were started from the outside to the state machines.
    -- * The InternalInvocationProxy processes dispatch invocations between state machines.

    -- Custom inter-dependent type declarations start
    type \unsigned32_Array\ is array (integer range <>) of unsigned(31 downto 0);
    type \Lombiq.Unum.BitMask\ is record 
        \IsNull\: boolean;
        \Size\: unsigned(15 downto 0);
        \SegmentCount\: unsigned(15 downto 0);
        \Segments\: \unsigned32_Array\(0 to 8);
    end record;
    type \Lombiq.Unum.UnumEnvironment\ is record 
        \IsNull\: boolean;
        \ExponentSizeSize\: unsigned(7 downto 0);
        \FractionSizeSize\: unsigned(7 downto 0);
        \ExponentSizeMax\: unsigned(7 downto 0);
        \FractionSizeMax\: unsigned(15 downto 0);
        \UnumTagSize\: unsigned(7 downto 0);
        \Size\: unsigned(15 downto 0);
        \EmptyBitMask\: \Lombiq.Unum.BitMask\;
        \UncertaintyBitMask\: \Lombiq.Unum.BitMask\;
        \ExponentSizeMask\: \Lombiq.Unum.BitMask\;
        \FractionSizeMask\: \Lombiq.Unum.BitMask\;
        \ExponentAndFractionSizeMask\: \Lombiq.Unum.BitMask\;
        \UnumTagMask\: \Lombiq.Unum.BitMask\;
        \SignBitMask\: \Lombiq.Unum.BitMask\;
        \ULP\: \Lombiq.Unum.BitMask\;
        \PositiveInfinity\: \Lombiq.Unum.BitMask\;
        \NegativeInfinity\: \Lombiq.Unum.BitMask\;
        \QuietNotANumber\: \Lombiq.Unum.BitMask\;
        \SignalingNotANumber\: \Lombiq.Unum.BitMask\;
        \LargestPositive\: \Lombiq.Unum.BitMask\;
        \SmallestPositive\: \Lombiq.Unum.BitMask\;
        \LargestNegative\: \Lombiq.Unum.BitMask\;
        \MinRealU\: \Lombiq.Unum.BitMask\;
    end record;
    type \Lombiq.Unum.Unum\ is record 
        \IsNull\: boolean;
        \_environment\: \Lombiq.Unum.UnumEnvironment\;
        \UnumBits\: \Lombiq.Unum.BitMask\;
    end record;
    -- Custom inter-dependent type declarations end


    -- System.Void Hast.Samples.SampleAssembly.UnumCalculator::CalculateSumOfPowersofTwo(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations start
    -- State machine states:
    type \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._States\ is (
        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_0\, 
        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_1\, 
        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_2\, 
        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_3\, 
        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_4\, 
        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_5\, 
        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_6\, 
        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_7\, 
        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_8\, 
        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_9\, 
        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_10\, 
        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_11\, 
        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_12\, 
        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_13\, 
        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_14\, 
        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_15\, 
        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_16\);
    -- Signals:
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._Finished\: boolean := false;
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.SimpleMemory.DataOut\: std_logic_vector(31 downto 0);
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.SimpleMemory.ReadEnable\: boolean := false;
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.SimpleMemory.WriteEnable\: boolean := false;
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.UnumCalculator::EnvironmentFactory()._Started.0\: boolean := false;
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32).this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32).environment.parameter.Out.0\: \Lombiq.Unum.UnumEnvironment\;
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32).value.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32)._Started.0\: boolean := false;
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum).left.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum).right.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum)._Started.0\: boolean := false;
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::FractionToUintArray().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::FractionToUintArray()._Started.0\: boolean := false;
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._Started\: boolean := false;
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.UnumCalculator::EnvironmentFactory()._Finished.0\: boolean := false;
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.UnumCalculator::EnvironmentFactory().return.0\: \Lombiq.Unum.UnumEnvironment\;
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32).this.parameter.In.0\: \Lombiq.Unum.Unum\;
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32).environment.parameter.In.0\: \Lombiq.Unum.UnumEnvironment\;
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32)._Finished.0\: boolean := false;
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum)._Finished.0\: boolean := false;
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum).return.0\: \Lombiq.Unum.Unum\;
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::FractionToUintArray()._Finished.0\: boolean := false;
    Signal \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::FractionToUintArray().return.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    -- System.Void Hast.Samples.SampleAssembly.UnumCalculator::CalculateSumOfPowersofTwo(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 declarations end


    -- Lombiq.Unum.UnumEnvironment Hast.Samples.SampleAssembly.UnumCalculator::EnvironmentFactory().0 declarations start
    -- State machine states:
    type \UnumCalculator::EnvironmentFactory().0._States\ is (
        \UnumCalculator::EnvironmentFactory().0._State_0\, 
        \UnumCalculator::EnvironmentFactory().0._State_1\, 
        \UnumCalculator::EnvironmentFactory().0._State_2\, 
        \UnumCalculator::EnvironmentFactory().0._State_3\);
    -- Signals:
    Signal \UnumCalculator::EnvironmentFactory().0._Finished\: boolean := false;
    Signal \UnumCalculator::EnvironmentFactory().0.return\: \Lombiq.Unum.UnumEnvironment\;
    Signal \UnumCalculator::EnvironmentFactory().0.UnumEnvironment::.ctor(Byte,Byte).this.parameter.Out.0\: \Lombiq.Unum.UnumEnvironment\;
    Signal \UnumCalculator::EnvironmentFactory().0.UnumEnvironment::.ctor(Byte,Byte).exponentSizeSize.parameter.Out.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
    Signal \UnumCalculator::EnvironmentFactory().0.UnumEnvironment::.ctor(Byte,Byte).fractionSizeSize.parameter.Out.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
    Signal \UnumCalculator::EnvironmentFactory().0.UnumEnvironment::.ctor(Byte,Byte)._Started.0\: boolean := false;
    Signal \UnumCalculator::EnvironmentFactory().0._Started\: boolean := false;
    Signal \UnumCalculator::EnvironmentFactory().0.UnumEnvironment::.ctor(Byte,Byte).this.parameter.In.0\: \Lombiq.Unum.UnumEnvironment\;
    Signal \UnumCalculator::EnvironmentFactory().0.UnumEnvironment::.ctor(Byte,Byte)._Finished.0\: boolean := false;
    -- Lombiq.Unum.UnumEnvironment Hast.Samples.SampleAssembly.UnumCalculator::EnvironmentFactory().0 declarations end


    -- System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16).0 declarations start
    -- State machine states:
    type \BitMask::.ctor(UInt32[],UInt16).0._States\ is (
        \BitMask::.ctor(UInt32[],UInt16).0._State_0\, 
        \BitMask::.ctor(UInt32[],UInt16).0._State_1\, 
        \BitMask::.ctor(UInt32[],UInt16).0._State_2\, 
        \BitMask::.ctor(UInt32[],UInt16).0._State_3\, 
        \BitMask::.ctor(UInt32[],UInt16).0._State_4\, 
        \BitMask::.ctor(UInt32[],UInt16).0._State_5\, 
        \BitMask::.ctor(UInt32[],UInt16).0._State_6\, 
        \BitMask::.ctor(UInt32[],UInt16).0._State_7\, 
        \BitMask::.ctor(UInt32[],UInt16).0._State_8\, 
        \BitMask::.ctor(UInt32[],UInt16).0._State_9\, 
        \BitMask::.ctor(UInt32[],UInt16).0._State_10\, 
        \BitMask::.ctor(UInt32[],UInt16).0._State_11\, 
        \BitMask::.ctor(UInt32[],UInt16).0._State_12\, 
        \BitMask::.ctor(UInt32[],UInt16).0._State_13\, 
        \BitMask::.ctor(UInt32[],UInt16).0._State_14\, 
        \BitMask::.ctor(UInt32[],UInt16).0._State_15\, 
        \BitMask::.ctor(UInt32[],UInt16).0._State_16\);
    -- Signals:
    Signal \BitMask::.ctor(UInt32[],UInt16).0._Finished\: boolean := false;
    Signal \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.Out\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.Out\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::.ctor(UInt32[],UInt16).0._Started\: boolean := false;
    Signal \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.In\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::.ctor(UInt32[],UInt16).0.size.parameter.In\: unsigned(15 downto 0) := to_unsigned(0, 16);
    -- System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16).0 declarations end


    -- System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean).0 declarations start
    -- State machine states:
    type \BitMask::.ctor(UInt16,Boolean).0._States\ is (
        \BitMask::.ctor(UInt16,Boolean).0._State_0\, 
        \BitMask::.ctor(UInt16,Boolean).0._State_1\, 
        \BitMask::.ctor(UInt16,Boolean).0._State_2\, 
        \BitMask::.ctor(UInt16,Boolean).0._State_3\, 
        \BitMask::.ctor(UInt16,Boolean).0._State_4\, 
        \BitMask::.ctor(UInt16,Boolean).0._State_5\, 
        \BitMask::.ctor(UInt16,Boolean).0._State_6\, 
        \BitMask::.ctor(UInt16,Boolean).0._State_7\);
    -- Signals:
    Signal \BitMask::.ctor(UInt16,Boolean).0._Finished\: boolean := false;
    Signal \BitMask::.ctor(UInt16,Boolean).0.this.parameter.Out\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::.ctor(UInt16,Boolean).0._Started\: boolean := false;
    Signal \BitMask::.ctor(UInt16,Boolean).0.this.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::.ctor(UInt16,Boolean).0.size.parameter.In\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \BitMask::.ctor(UInt16,Boolean).0.allOne.parameter.In\: boolean := false;
    -- System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean).0 declarations end


    -- System.Void Lombiq.Unum.BitMask::.ctor(Lombiq.Unum.BitMask).0 declarations start
    -- State machine states:
    type \BitMask::.ctor(BitMask).0._States\ is (
        \BitMask::.ctor(BitMask).0._State_0\, 
        \BitMask::.ctor(BitMask).0._State_1\, 
        \BitMask::.ctor(BitMask).0._State_2\);
    -- Signals:
    Signal \BitMask::.ctor(BitMask).0._Finished\: boolean := false;
    Signal \BitMask::.ctor(BitMask).0.this.parameter.Out\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::.ctor(BitMask).0.source.parameter.Out\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::.ctor(BitMask).0._Started\: boolean := false;
    Signal \BitMask::.ctor(BitMask).0.this.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::.ctor(BitMask).0.source.parameter.In\: \Lombiq.Unum.BitMask\;
    -- System.Void Lombiq.Unum.BitMask::.ctor(Lombiq.Unum.BitMask).0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::FromImmutableArray(System.UInt32[],System.UInt16).0 declarations start
    -- State machine states:
    type \BitMask::FromImmutableArray(UInt32[],UInt16).0._States\ is (
        \BitMask::FromImmutableArray(UInt32[],UInt16).0._State_0\, 
        \BitMask::FromImmutableArray(UInt32[],UInt16).0._State_1\, 
        \BitMask::FromImmutableArray(UInt32[],UInt16).0._State_2\, 
        \BitMask::FromImmutableArray(UInt32[],UInt16).0._State_3\);
    -- Signals:
    Signal \BitMask::FromImmutableArray(UInt32[],UInt16).0._Finished\: boolean := false;
    Signal \BitMask::FromImmutableArray(UInt32[],UInt16).0.return\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::FromImmutableArray(UInt32[],UInt16).0.segments.parameter.Out\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\: boolean := false;
    Signal \BitMask::FromImmutableArray(UInt32[],UInt16).0._Started\: boolean := false;
    Signal \BitMask::FromImmutableArray(UInt32[],UInt16).0.segments.parameter.In\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::FromImmutableArray(UInt32[],UInt16).0.size.parameter.In\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\: boolean := false;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::FromImmutableArray(System.UInt32[],System.UInt16).0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetOne(System.UInt16).0 declarations start
    -- State machine states:
    type \BitMask::SetOne(UInt16).0._States\ is (
        \BitMask::SetOne(UInt16).0._State_0\, 
        \BitMask::SetOne(UInt16).0._State_1\, 
        \BitMask::SetOne(UInt16).0._State_2\, 
        \BitMask::SetOne(UInt16).0._State_3\, 
        \BitMask::SetOne(UInt16).0._State_4\, 
        \BitMask::SetOne(UInt16).0._State_5\, 
        \BitMask::SetOne(UInt16).0._State_6\, 
        \BitMask::SetOne(UInt16).0._State_7\, 
        \BitMask::SetOne(UInt16).0._State_8\, 
        \BitMask::SetOne(UInt16).0._State_9\, 
        \BitMask::SetOne(UInt16).0._State_10\, 
        \BitMask::SetOne(UInt16).0._State_11\, 
        \BitMask::SetOne(UInt16).0._State_12\, 
        \BitMask::SetOne(UInt16).0._State_13\, 
        \BitMask::SetOne(UInt16).0._State_14\, 
        \BitMask::SetOne(UInt16).0._State_15\);
    -- Signals:
    Signal \BitMask::SetOne(UInt16).0._Finished\: boolean := false;
    Signal \BitMask::SetOne(UInt16).0.return\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask).source.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask)._Started.0\: boolean := false;
    Signal \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).segments.parameter.Out.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Started.0\: boolean := false;
    Signal \BitMask::SetOne(UInt16).0._Started\: boolean := false;
    Signal \BitMask::SetOne(UInt16).0.this.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::SetOne(UInt16).0.index.parameter.In\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask).this.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask).source.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask)._Finished.0\: boolean := false;
    Signal \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).segments.parameter.In.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Finished.0\: boolean := false;
    Signal \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).return.0\: \Lombiq.Unum.BitMask\;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetOne(System.UInt16).0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetZero(System.UInt16).0 declarations start
    -- State machine states:
    type \BitMask::SetZero(UInt16).0._States\ is (
        \BitMask::SetZero(UInt16).0._State_0\, 
        \BitMask::SetZero(UInt16).0._State_1\, 
        \BitMask::SetZero(UInt16).0._State_2\, 
        \BitMask::SetZero(UInt16).0._State_3\, 
        \BitMask::SetZero(UInt16).0._State_4\, 
        \BitMask::SetZero(UInt16).0._State_5\, 
        \BitMask::SetZero(UInt16).0._State_6\, 
        \BitMask::SetZero(UInt16).0._State_7\, 
        \BitMask::SetZero(UInt16).0._State_8\, 
        \BitMask::SetZero(UInt16).0._State_9\, 
        \BitMask::SetZero(UInt16).0._State_10\, 
        \BitMask::SetZero(UInt16).0._State_11\, 
        \BitMask::SetZero(UInt16).0._State_12\, 
        \BitMask::SetZero(UInt16).0._State_13\, 
        \BitMask::SetZero(UInt16).0._State_14\, 
        \BitMask::SetZero(UInt16).0._State_15\);
    -- Signals:
    Signal \BitMask::SetZero(UInt16).0._Finished\: boolean := false;
    Signal \BitMask::SetZero(UInt16).0.return\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask).source.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask)._Started.0\: boolean := false;
    Signal \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).segments.parameter.Out.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Started.0\: boolean := false;
    Signal \BitMask::SetZero(UInt16).0._Started\: boolean := false;
    Signal \BitMask::SetZero(UInt16).0.this.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::SetZero(UInt16).0.index.parameter.In\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask).this.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask).source.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask)._Finished.0\: boolean := false;
    Signal \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).segments.parameter.In.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Finished.0\: boolean := false;
    Signal \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).return.0\: \Lombiq.Unum.BitMask\;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetZero(System.UInt16).0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::ShiftOutLeastSignificantZeros().0 declarations start
    -- State machine states:
    type \BitMask::ShiftOutLeastSignificantZeros().0._States\ is (
        \BitMask::ShiftOutLeastSignificantZeros().0._State_0\, 
        \BitMask::ShiftOutLeastSignificantZeros().0._State_1\, 
        \BitMask::ShiftOutLeastSignificantZeros().0._State_2\, 
        \BitMask::ShiftOutLeastSignificantZeros().0._State_3\, 
        \BitMask::ShiftOutLeastSignificantZeros().0._State_4\, 
        \BitMask::ShiftOutLeastSignificantZeros().0._State_5\, 
        \BitMask::ShiftOutLeastSignificantZeros().0._State_6\, 
        \BitMask::ShiftOutLeastSignificantZeros().0._State_7\, 
        \BitMask::ShiftOutLeastSignificantZeros().0._State_8\);
    -- Signals:
    Signal \BitMask::ShiftOutLeastSignificantZeros().0._Finished\: boolean := false;
    Signal \BitMask::ShiftOutLeastSignificantZeros().0.return\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::GetLeastSignificantOnePosition().this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::GetLeastSignificantOnePosition()._Started.0\: boolean := false;
    Signal \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask).source.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask)._Started.0\: boolean := false;
    Signal \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::op_RightShift(BitMask,Int32).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::op_RightShift(BitMask,Int32).right.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\: boolean := false;
    Signal \BitMask::ShiftOutLeastSignificantZeros().0._Started\: boolean := false;
    Signal \BitMask::ShiftOutLeastSignificantZeros().0.this.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::GetLeastSignificantOnePosition()._Finished.0\: boolean := false;
    Signal \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::GetLeastSignificantOnePosition().return.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask).this.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask).source.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask)._Finished.0\: boolean := false;
    Signal \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\: boolean := false;
    Signal \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::op_RightShift(BitMask,Int32).return.0\: \Lombiq.Unum.BitMask\;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::ShiftOutLeastSignificantZeros().0 declarations end


    -- System.Boolean Lombiq.Unum.BitMask::op_Equality(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 declarations start
    -- State machine states:
    type \BitMask::op_Equality(BitMask,BitMask).0._States\ is (
        \BitMask::op_Equality(BitMask,BitMask).0._State_0\, 
        \BitMask::op_Equality(BitMask,BitMask).0._State_1\, 
        \BitMask::op_Equality(BitMask,BitMask).0._State_2\, 
        \BitMask::op_Equality(BitMask,BitMask).0._State_3\, 
        \BitMask::op_Equality(BitMask,BitMask).0._State_4\, 
        \BitMask::op_Equality(BitMask,BitMask).0._State_5\, 
        \BitMask::op_Equality(BitMask,BitMask).0._State_6\, 
        \BitMask::op_Equality(BitMask,BitMask).0._State_7\, 
        \BitMask::op_Equality(BitMask,BitMask).0._State_8\, 
        \BitMask::op_Equality(BitMask,BitMask).0._State_9\);
    -- Signals:
    Signal \BitMask::op_Equality(BitMask,BitMask).0._Finished\: boolean := false;
    Signal \BitMask::op_Equality(BitMask,BitMask).0.return\: boolean := false;
    Signal \BitMask::op_Equality(BitMask,BitMask).0._Started\: boolean := false;
    Signal \BitMask::op_Equality(BitMask,BitMask).0.left.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_Equality(BitMask,BitMask).0.right.parameter.In\: \Lombiq.Unum.BitMask\;
    -- System.Boolean Lombiq.Unum.BitMask::op_Equality(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 declarations end


    -- System.Boolean Lombiq.Unum.BitMask::op_GreaterThan(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 declarations start
    -- State machine states:
    type \BitMask::op_GreaterThan(BitMask,BitMask).0._States\ is (
        \BitMask::op_GreaterThan(BitMask,BitMask).0._State_0\, 
        \BitMask::op_GreaterThan(BitMask,BitMask).0._State_1\, 
        \BitMask::op_GreaterThan(BitMask,BitMask).0._State_2\, 
        \BitMask::op_GreaterThan(BitMask,BitMask).0._State_3\, 
        \BitMask::op_GreaterThan(BitMask,BitMask).0._State_4\, 
        \BitMask::op_GreaterThan(BitMask,BitMask).0._State_5\, 
        \BitMask::op_GreaterThan(BitMask,BitMask).0._State_6\);
    -- Signals:
    Signal \BitMask::op_GreaterThan(BitMask,BitMask).0._Finished\: boolean := false;
    Signal \BitMask::op_GreaterThan(BitMask,BitMask).0.return\: boolean := false;
    Signal \BitMask::op_GreaterThan(BitMask,BitMask).0._Started\: boolean := false;
    Signal \BitMask::op_GreaterThan(BitMask,BitMask).0.left.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_GreaterThan(BitMask,BitMask).0.right.parameter.In\: \Lombiq.Unum.BitMask\;
    -- System.Boolean Lombiq.Unum.BitMask::op_GreaterThan(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 declarations end


    -- System.Boolean Lombiq.Unum.BitMask::op_LessThan(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 declarations start
    -- State machine states:
    type \BitMask::op_LessThan(BitMask,BitMask).0._States\ is (
        \BitMask::op_LessThan(BitMask,BitMask).0._State_0\, 
        \BitMask::op_LessThan(BitMask,BitMask).0._State_1\, 
        \BitMask::op_LessThan(BitMask,BitMask).0._State_2\, 
        \BitMask::op_LessThan(BitMask,BitMask).0._State_3\, 
        \BitMask::op_LessThan(BitMask,BitMask).0._State_4\, 
        \BitMask::op_LessThan(BitMask,BitMask).0._State_5\, 
        \BitMask::op_LessThan(BitMask,BitMask).0._State_6\);
    -- Signals:
    Signal \BitMask::op_LessThan(BitMask,BitMask).0._Finished\: boolean := false;
    Signal \BitMask::op_LessThan(BitMask,BitMask).0.return\: boolean := false;
    Signal \BitMask::op_LessThan(BitMask,BitMask).0._Started\: boolean := false;
    Signal \BitMask::op_LessThan(BitMask,BitMask).0.left.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_LessThan(BitMask,BitMask).0.right.parameter.In\: \Lombiq.Unum.BitMask\;
    -- System.Boolean Lombiq.Unum.BitMask::op_LessThan(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 declarations end


    -- System.Boolean Lombiq.Unum.BitMask::op_GreaterThanOrEqual(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 declarations start
    -- State machine states:
    type \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._States\ is (
        \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._State_0\, 
        \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._State_1\, 
        \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._State_2\, 
        \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._State_3\);
    -- Signals:
    Signal \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._Finished\: boolean := false;
    Signal \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.return\: boolean := false;
    Signal \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.BitMask::op_LessThan(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.BitMask::op_LessThan(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.BitMask::op_LessThan(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._Started\: boolean := false;
    Signal \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.left.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.right.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.BitMask::op_LessThan(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.BitMask::op_LessThan(BitMask,BitMask).return.0\: boolean := false;
    -- System.Boolean Lombiq.Unum.BitMask::op_GreaterThanOrEqual(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,System.UInt32).0 declarations start
    -- State machine states:
    type \BitMask::op_Addition(BitMask,UInt32).0._States\ is (
        \BitMask::op_Addition(BitMask,UInt32).0._State_0\, 
        \BitMask::op_Addition(BitMask,UInt32).0._State_1\, 
        \BitMask::op_Addition(BitMask,UInt32).0._State_2\, 
        \BitMask::op_Addition(BitMask,UInt32).0._State_3\, 
        \BitMask::op_Addition(BitMask,UInt32).0._State_4\);
    -- Signals:
    Signal \BitMask::op_Addition(BitMask,UInt32).0._Finished\: boolean := false;
    Signal \BitMask::op_Addition(BitMask,UInt32).0.return\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\: boolean := false;
    Signal \BitMask::op_Addition(BitMask,UInt32).0.BitMask::op_Addition(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_Addition(BitMask,UInt32).0.BitMask::op_Addition(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_Addition(BitMask,UInt32).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \BitMask::op_Addition(BitMask,UInt32).0._Started\: boolean := false;
    Signal \BitMask::op_Addition(BitMask,UInt32).0.left.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_Addition(BitMask,UInt32).0.right.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\: boolean := false;
    Signal \BitMask::op_Addition(BitMask,UInt32).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \BitMask::op_Addition(BitMask,UInt32).0.BitMask::op_Addition(BitMask,BitMask).return.0\: \Lombiq.Unum.BitMask\;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,System.UInt32).0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,System.UInt32).0 declarations start
    -- State machine states:
    type \BitMask::op_Subtraction(BitMask,UInt32).0._States\ is (
        \BitMask::op_Subtraction(BitMask,UInt32).0._State_0\, 
        \BitMask::op_Subtraction(BitMask,UInt32).0._State_1\, 
        \BitMask::op_Subtraction(BitMask,UInt32).0._State_2\, 
        \BitMask::op_Subtraction(BitMask,UInt32).0._State_3\, 
        \BitMask::op_Subtraction(BitMask,UInt32).0._State_4\);
    -- Signals:
    Signal \BitMask::op_Subtraction(BitMask,UInt32).0._Finished\: boolean := false;
    Signal \BitMask::op_Subtraction(BitMask,UInt32).0.return\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\: boolean := false;
    Signal \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::op_Subtraction(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::op_Subtraction(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \BitMask::op_Subtraction(BitMask,UInt32).0._Started\: boolean := false;
    Signal \BitMask::op_Subtraction(BitMask,UInt32).0.left.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_Subtraction(BitMask,UInt32).0.right.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\: boolean := false;
    Signal \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::op_Subtraction(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::op_Subtraction(BitMask,BitMask).return.0\: \Lombiq.Unum.BitMask\;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,System.UInt32).0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 declarations start
    -- State machine states:
    type \BitMask::op_Addition(BitMask,BitMask).0._States\ is (
        \BitMask::op_Addition(BitMask,BitMask).0._State_0\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_1\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_2\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_3\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_4\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_5\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_6\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_7\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_8\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_9\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_10\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_11\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_12\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_13\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_14\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_15\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_16\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_17\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_18\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_19\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_20\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_21\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_22\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_23\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_24\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_25\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_26\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_27\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_28\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_29\, 
        \BitMask::op_Addition(BitMask,BitMask).0._State_30\);
    -- Signals:
    Signal \BitMask::op_Addition(BitMask,BitMask).0._Finished\: boolean := false;
    Signal \BitMask::op_Addition(BitMask,BitMask).0.return\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\: boolean := false;
    Signal \BitMask::op_Addition(BitMask,BitMask).0._Started\: boolean := false;
    Signal \BitMask::op_Addition(BitMask,BitMask).0.left.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_Addition(BitMask,BitMask).0.right.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\: boolean := false;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 declarations start
    -- State machine states:
    type \BitMask::op_Subtraction(BitMask,BitMask).0._States\ is (
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_0\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_1\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_2\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_3\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_4\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_5\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_6\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_7\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_8\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_9\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_10\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_11\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_12\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_13\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_14\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_15\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_16\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_17\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_18\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_19\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_20\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_21\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_22\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_23\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_24\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_25\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_26\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_27\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_28\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_29\, 
        \BitMask::op_Subtraction(BitMask,BitMask).0._State_30\);
    -- Signals:
    Signal \BitMask::op_Subtraction(BitMask,BitMask).0._Finished\: boolean := false;
    Signal \BitMask::op_Subtraction(BitMask,BitMask).0.return\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\: boolean := false;
    Signal \BitMask::op_Subtraction(BitMask,BitMask).0._Started\: boolean := false;
    Signal \BitMask::op_Subtraction(BitMask,BitMask).0.left.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_Subtraction(BitMask,BitMask).0.right.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\: boolean := false;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseOr(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 declarations start
    -- State machine states:
    type \BitMask::op_BitwiseOr(BitMask,BitMask).0._States\ is (
        \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_0\, 
        \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_1\, 
        \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_2\, 
        \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_3\, 
        \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_4\, 
        \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_5\, 
        \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_6\, 
        \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_7\, 
        \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_8\, 
        \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_9\);
    -- Signals:
    Signal \BitMask::op_BitwiseOr(BitMask,BitMask).0._Finished\: boolean := false;
    Signal \BitMask::op_BitwiseOr(BitMask,BitMask).0.return\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\: boolean := false;
    Signal \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Started.0\: boolean := false;
    Signal \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\: boolean := false;
    Signal \BitMask::op_BitwiseOr(BitMask,BitMask).0._Started\: boolean := false;
    Signal \BitMask::op_BitwiseOr(BitMask,BitMask).0.left.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_BitwiseOr(BitMask,BitMask).0.right.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\: boolean := false;
    Signal \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\: boolean := false;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseOr(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseAnd(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 declarations start
    -- State machine states:
    type \BitMask::op_BitwiseAnd(BitMask,BitMask).0._States\ is (
        \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_0\, 
        \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_1\, 
        \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_2\, 
        \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_3\, 
        \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_4\, 
        \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_5\, 
        \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_6\, 
        \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_7\, 
        \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_8\, 
        \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_9\);
    -- Signals:
    Signal \BitMask::op_BitwiseAnd(BitMask,BitMask).0._Finished\: boolean := false;
    Signal \BitMask::op_BitwiseAnd(BitMask,BitMask).0.return\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\: boolean := false;
    Signal \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Started.0\: boolean := false;
    Signal \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\: boolean := false;
    Signal \BitMask::op_BitwiseAnd(BitMask,BitMask).0._Started\: boolean := false;
    Signal \BitMask::op_BitwiseAnd(BitMask,BitMask).0.left.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_BitwiseAnd(BitMask,BitMask).0.right.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\: boolean := false;
    Signal \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\: boolean := false;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseAnd(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_RightShift(Lombiq.Unum.BitMask,System.Int32).0 declarations start
    -- State machine states:
    type \BitMask::op_RightShift(BitMask,Int32).0._States\ is (
        \BitMask::op_RightShift(BitMask,Int32).0._State_0\, 
        \BitMask::op_RightShift(BitMask,Int32).0._State_1\, 
        \BitMask::op_RightShift(BitMask,Int32).0._State_2\, 
        \BitMask::op_RightShift(BitMask,Int32).0._State_3\, 
        \BitMask::op_RightShift(BitMask,Int32).0._State_4\, 
        \BitMask::op_RightShift(BitMask,Int32).0._State_5\, 
        \BitMask::op_RightShift(BitMask,Int32).0._State_6\, 
        \BitMask::op_RightShift(BitMask,Int32).0._State_7\, 
        \BitMask::op_RightShift(BitMask,Int32).0._State_8\, 
        \BitMask::op_RightShift(BitMask,Int32).0._State_9\, 
        \BitMask::op_RightShift(BitMask,Int32).0._State_10\, 
        \BitMask::op_RightShift(BitMask,Int32).0._State_11\, 
        \BitMask::op_RightShift(BitMask,Int32).0._State_12\, 
        \BitMask::op_RightShift(BitMask,Int32).0._State_13\, 
        \BitMask::op_RightShift(BitMask,Int32).0._State_14\, 
        \BitMask::op_RightShift(BitMask,Int32).0._State_15\);
    -- Signals:
    Signal \BitMask::op_RightShift(BitMask,Int32).0._Finished\: boolean := false;
    Signal \BitMask::op_RightShift(BitMask,Int32).0.return\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_RightShift(BitMask,Int32).0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_RightShift(BitMask,Int32).0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \BitMask::op_RightShift(BitMask,Int32).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\: boolean := false;
    Signal \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\: boolean := false;
    Signal \BitMask::op_RightShift(BitMask,Int32).0._Started\: boolean := false;
    Signal \BitMask::op_RightShift(BitMask,Int32).0.left.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_RightShift(BitMask,Int32).0.right.parameter.In\: signed(31 downto 0) := to_signed(0, 32);
    Signal \BitMask::op_RightShift(BitMask,Int32).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\: boolean := false;
    Signal \BitMask::op_RightShift(BitMask,Int32).0.BitMask::op_LeftShift(BitMask,Int32).return.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\: boolean := false;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_RightShift(Lombiq.Unum.BitMask,System.Int32).0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32).0 declarations start
    -- State machine states:
    type \BitMask::op_LeftShift(BitMask,Int32).0._States\ is (
        \BitMask::op_LeftShift(BitMask,Int32).0._State_0\, 
        \BitMask::op_LeftShift(BitMask,Int32).0._State_1\, 
        \BitMask::op_LeftShift(BitMask,Int32).0._State_2\, 
        \BitMask::op_LeftShift(BitMask,Int32).0._State_3\, 
        \BitMask::op_LeftShift(BitMask,Int32).0._State_4\, 
        \BitMask::op_LeftShift(BitMask,Int32).0._State_5\, 
        \BitMask::op_LeftShift(BitMask,Int32).0._State_6\, 
        \BitMask::op_LeftShift(BitMask,Int32).0._State_7\, 
        \BitMask::op_LeftShift(BitMask,Int32).0._State_8\, 
        \BitMask::op_LeftShift(BitMask,Int32).0._State_9\, 
        \BitMask::op_LeftShift(BitMask,Int32).0._State_10\, 
        \BitMask::op_LeftShift(BitMask,Int32).0._State_11\, 
        \BitMask::op_LeftShift(BitMask,Int32).0._State_12\, 
        \BitMask::op_LeftShift(BitMask,Int32).0._State_13\);
    -- Signals:
    Signal \BitMask::op_LeftShift(BitMask,Int32).0._Finished\: boolean := false;
    Signal \BitMask::op_LeftShift(BitMask,Int32).0.return\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::op_RightShift(BitMask,Int32).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::op_RightShift(BitMask,Int32).right.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::op_RightShift(BitMask,Int32)._Started.0\: boolean := false;
    Signal \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\: boolean := false;
    Signal \BitMask::op_LeftShift(BitMask,Int32).0._Started\: boolean := false;
    Signal \BitMask::op_LeftShift(BitMask,Int32).0.left.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_LeftShift(BitMask,Int32).0.right.parameter.In\: signed(31 downto 0) := to_signed(0, 32);
    Signal \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\: boolean := false;
    Signal \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::op_RightShift(BitMask,Int32).return.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\: boolean := false;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32).0 declarations end


    -- System.UInt16 Lombiq.Unum.BitMask::GetMostSignificantOnePosition().0 declarations start
    -- State machine states:
    type \BitMask::GetMostSignificantOnePosition().0._States\ is (
        \BitMask::GetMostSignificantOnePosition().0._State_0\, 
        \BitMask::GetMostSignificantOnePosition().0._State_1\, 
        \BitMask::GetMostSignificantOnePosition().0._State_2\, 
        \BitMask::GetMostSignificantOnePosition().0._State_3\, 
        \BitMask::GetMostSignificantOnePosition().0._State_4\, 
        \BitMask::GetMostSignificantOnePosition().0._State_5\, 
        \BitMask::GetMostSignificantOnePosition().0._State_6\, 
        \BitMask::GetMostSignificantOnePosition().0._State_7\, 
        \BitMask::GetMostSignificantOnePosition().0._State_8\);
    -- Signals:
    Signal \BitMask::GetMostSignificantOnePosition().0._Finished\: boolean := false;
    Signal \BitMask::GetMostSignificantOnePosition().0.return\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \BitMask::GetMostSignificantOnePosition().0._Started\: boolean := false;
    Signal \BitMask::GetMostSignificantOnePosition().0.this.parameter.In\: \Lombiq.Unum.BitMask\;
    -- System.UInt16 Lombiq.Unum.BitMask::GetMostSignificantOnePosition().0 declarations end


    -- System.UInt16 Lombiq.Unum.BitMask::GetLeastSignificantOnePosition().0 declarations start
    -- State machine states:
    type \BitMask::GetLeastSignificantOnePosition().0._States\ is (
        \BitMask::GetLeastSignificantOnePosition().0._State_0\, 
        \BitMask::GetLeastSignificantOnePosition().0._State_1\, 
        \BitMask::GetLeastSignificantOnePosition().0._State_2\, 
        \BitMask::GetLeastSignificantOnePosition().0._State_3\, 
        \BitMask::GetLeastSignificantOnePosition().0._State_4\, 
        \BitMask::GetLeastSignificantOnePosition().0._State_5\, 
        \BitMask::GetLeastSignificantOnePosition().0._State_6\, 
        \BitMask::GetLeastSignificantOnePosition().0._State_7\, 
        \BitMask::GetLeastSignificantOnePosition().0._State_8\, 
        \BitMask::GetLeastSignificantOnePosition().0._State_9\, 
        \BitMask::GetLeastSignificantOnePosition().0._State_10\, 
        \BitMask::GetLeastSignificantOnePosition().0._State_11\, 
        \BitMask::GetLeastSignificantOnePosition().0._State_12\, 
        \BitMask::GetLeastSignificantOnePosition().0._State_13\, 
        \BitMask::GetLeastSignificantOnePosition().0._State_14\, 
        \BitMask::GetLeastSignificantOnePosition().0._State_15\, 
        \BitMask::GetLeastSignificantOnePosition().0._State_16\, 
        \BitMask::GetLeastSignificantOnePosition().0._State_17\);
    -- Signals:
    Signal \BitMask::GetLeastSignificantOnePosition().0._Finished\: boolean := false;
    Signal \BitMask::GetLeastSignificantOnePosition().0.return\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \BitMask::GetLeastSignificantOnePosition().0._Started\: boolean := false;
    Signal \BitMask::GetLeastSignificantOnePosition().0.this.parameter.In\: \Lombiq.Unum.BitMask\;
    -- System.UInt16 Lombiq.Unum.BitMask::GetLeastSignificantOnePosition().0 declarations end


    -- System.UInt32 Lombiq.Unum.BitMask::GetLowest32Bits().0 declarations start
    -- State machine states:
    type \BitMask::GetLowest32Bits().0._States\ is (
        \BitMask::GetLowest32Bits().0._State_0\, 
        \BitMask::GetLowest32Bits().0._State_1\, 
        \BitMask::GetLowest32Bits().0._State_2\);
    -- Signals:
    Signal \BitMask::GetLowest32Bits().0._Finished\: boolean := false;
    Signal \BitMask::GetLowest32Bits().0.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \BitMask::GetLowest32Bits().0._Started\: boolean := false;
    Signal \BitMask::GetLowest32Bits().0.this.parameter.In\: \Lombiq.Unum.BitMask\;
    -- System.UInt32 Lombiq.Unum.BitMask::GetLowest32Bits().0 declarations end


    -- System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment).0 declarations start
    -- State machine states:
    type \Unum::.ctor(UnumEnvironment).0._States\ is (
        \Unum::.ctor(UnumEnvironment).0._State_0\, 
        \Unum::.ctor(UnumEnvironment).0._State_1\, 
        \Unum::.ctor(UnumEnvironment).0._State_2\, 
        \Unum::.ctor(UnumEnvironment).0._State_3\);
    -- Signals:
    Signal \Unum::.ctor(UnumEnvironment).0._Finished\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment).0.this.parameter.Out\: \Lombiq.Unum.Unum\;
    Signal \Unum::.ctor(UnumEnvironment).0.environment.parameter.Out\: \Lombiq.Unum.UnumEnvironment\;
    Signal \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean)._Started.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment).0._Started\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment).0.this.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::.ctor(UnumEnvironment).0.environment.parameter.In\: \Lombiq.Unum.UnumEnvironment\;
    Signal \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\: boolean := false;
    -- System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment).0 declarations end


    -- System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,Lombiq.Unum.BitMask).0 declarations start
    -- State machine states:
    type \Unum::.ctor(UnumEnvironment,BitMask).0._States\ is (
        \Unum::.ctor(UnumEnvironment,BitMask).0._State_0\, 
        \Unum::.ctor(UnumEnvironment,BitMask).0._State_1\, 
        \Unum::.ctor(UnumEnvironment,BitMask).0._State_2\, 
        \Unum::.ctor(UnumEnvironment,BitMask).0._State_3\);
    -- Signals:
    Signal \Unum::.ctor(UnumEnvironment,BitMask).0._Finished\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,BitMask).0.this.parameter.Out\: \Lombiq.Unum.Unum\;
    Signal \Unum::.ctor(UnumEnvironment,BitMask).0.environment.parameter.Out\: \Lombiq.Unum.UnumEnvironment\;
    Signal \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16).segments.parameter.Out.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Started.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,BitMask).0._Started\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,BitMask).0.this.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::.ctor(UnumEnvironment,BitMask).0.environment.parameter.In\: \Lombiq.Unum.UnumEnvironment\;
    Signal \Unum::.ctor(UnumEnvironment,BitMask).0.bits.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16).segments.parameter.In.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Finished.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16).return.0\: \Lombiq.Unum.BitMask\;
    -- System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,Lombiq.Unum.BitMask).0 declarations end


    -- System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.UInt32[],System.Boolean).0 declarations start
    -- State machine states:
    type \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._States\ is (
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_0\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_1\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_2\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_3\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_4\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_5\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_6\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_7\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_8\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_9\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_10\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_11\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_12\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_13\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_14\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_15\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_16\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_17\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_18\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_19\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_20\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_21\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_22\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_23\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_24\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_25\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_26\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_27\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_28\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_29\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_30\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_31\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_32\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_33\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_34\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_35\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_36\, 
        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_37\);
    -- Signals:
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._Finished\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.this.parameter.Out\: \Lombiq.Unum.Unum\;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.environment.parameter.Out\: \Lombiq.Unum.UnumEnvironment\;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.value.parameter.Out\: \unsigned32_Array\(0 to 0) := (others => to_unsigned(0, 32));
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Equality(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Equality(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Equality(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size()._Started.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition().this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition()._Started.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits().this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits()._Started.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Addition(BitMask,UInt32).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::ShiftOutLeastSignificantZeros().this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::ShiftOutLeastSignificantZeros()._Started.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::SetZero(UInt16).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::SetZero(UInt16).index.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::SetZero(UInt16)._Started.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).signBit.parameter.Out.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).exponent.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).fraction.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).uncertainityBit.parameter.Out.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).exponentSize.parameter.Out.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).fractionSize.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Started.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._Started\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.this.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.environment.parameter.In\: \Lombiq.Unum.UnumEnvironment\;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.value.parameter.In\: \unsigned32_Array\(0 to 0) := (others => to_unsigned(0, 32));
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.negative.parameter.In\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Equality(BitMask,BitMask).return.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size()._Finished.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size().return.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition()._Finished.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition().return.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits()._Finished.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits().return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Addition(BitMask,UInt32).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::ShiftOutLeastSignificantZeros()._Finished.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::ShiftOutLeastSignificantZeros().return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::SetZero(UInt16)._Finished.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::SetZero(UInt16).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Finished.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).return.0\: \Lombiq.Unum.BitMask\;
    -- System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.UInt32[],System.Boolean).0 declarations end


    -- System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.Int32).0 declarations start
    -- State machine states:
    type \Unum::.ctor(UnumEnvironment,Int32).0._States\ is (
        \Unum::.ctor(UnumEnvironment,Int32).0._State_0\, 
        \Unum::.ctor(UnumEnvironment,Int32).0._State_1\, 
        \Unum::.ctor(UnumEnvironment,Int32).0._State_2\, 
        \Unum::.ctor(UnumEnvironment,Int32).0._State_3\, 
        \Unum::.ctor(UnumEnvironment,Int32).0._State_4\, 
        \Unum::.ctor(UnumEnvironment,Int32).0._State_5\, 
        \Unum::.ctor(UnumEnvironment,Int32).0._State_6\, 
        \Unum::.ctor(UnumEnvironment,Int32).0._State_7\);
    -- Signals:
    Signal \Unum::.ctor(UnumEnvironment,Int32).0._Finished\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,Int32).0.this.parameter.Out\: \Lombiq.Unum.Unum\;
    Signal \Unum::.ctor(UnumEnvironment,Int32).0.environment.parameter.Out\: \Lombiq.Unum.UnumEnvironment\;
    Signal \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).environment.parameter.Out.0\: \Lombiq.Unum.UnumEnvironment\;
    Signal \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).value.parameter.Out.0\: \unsigned32_Array\(0 to 0) := (others => to_unsigned(0, 32));
    Signal \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).negative.parameter.Out.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean)._Started.0\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,Int32).0._Started\: boolean := false;
    Signal \Unum::.ctor(UnumEnvironment,Int32).0.this.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::.ctor(UnumEnvironment,Int32).0.environment.parameter.In\: \Lombiq.Unum.UnumEnvironment\;
    Signal \Unum::.ctor(UnumEnvironment,Int32).0.value.parameter.In\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).this.parameter.In.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).environment.parameter.In.0\: \Lombiq.Unum.UnumEnvironment\;
    Signal \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).value.parameter.In.0\: \unsigned32_Array\(0 to 0) := (others => to_unsigned(0, 32));
    Signal \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean)._Finished.0\: boolean := false;
    -- System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.Int32).0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::SetUnumBits(System.Boolean,Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean,System.Byte,System.UInt16).0 declarations start
    -- State machine states:
    type \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._States\ is (
        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_0\, 
        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_1\, 
        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_2\, 
        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_3\, 
        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_4\, 
        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_5\, 
        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_6\, 
        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_7\, 
        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_8\, 
        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_9\, 
        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_10\, 
        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_11\, 
        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_12\, 
        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_13\, 
        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_14\, 
        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_15\, 
        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_16\, 
        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_17\, 
        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_18\, 
        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_19\, 
        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_20\);
    -- Signals:
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._Finished\: boolean := false;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return\: \Lombiq.Unum.BitMask\;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_Size().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_Size()._Started.0\: boolean := false;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\: boolean := false;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\: boolean := false;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,UInt32).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\: boolean := false;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_UncertaintyBitMask().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_UncertaintyBitMask()._Started.0\: boolean := false;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_SignBitMask().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_SignBitMask()._Started.0\: boolean := false;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._Started\: boolean := false;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.this.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.signBit.parameter.In\: boolean := false;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.exponent.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.fraction.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.uncertainityBit.parameter.In\: boolean := false;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.exponentSize.parameter.In\: unsigned(7 downto 0) := to_unsigned(0, 8);
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.fractionSize.parameter.In\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_Size()._Finished.0\: boolean := false;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_Size().return.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\: boolean := false;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\: boolean := false;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\: boolean := false;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,UInt32).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_UncertaintyBitMask()._Finished.0\: boolean := false;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_UncertaintyBitMask().return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_SignBitMask()._Finished.0\: boolean := false;
    Signal \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_SignBitMask().return.0\: \Lombiq.Unum.BitMask\;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::SetUnumBits(System.Boolean,Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean,System.Byte,System.UInt16).0 declarations end


    -- System.UInt32[] Lombiq.Unum.Unum::FractionToUintArray().0 declarations start
    -- State machine states:
    type \Unum::FractionToUintArray().0._States\ is (
        \Unum::FractionToUintArray().0._State_0\, 
        \Unum::FractionToUintArray().0._State_1\, 
        \Unum::FractionToUintArray().0._State_2\, 
        \Unum::FractionToUintArray().0._State_3\, 
        \Unum::FractionToUintArray().0._State_4\, 
        \Unum::FractionToUintArray().0._State_5\, 
        \Unum::FractionToUintArray().0._State_6\, 
        \Unum::FractionToUintArray().0._State_7\, 
        \Unum::FractionToUintArray().0._State_8\, 
        \Unum::FractionToUintArray().0._State_9\, 
        \Unum::FractionToUintArray().0._State_10\, 
        \Unum::FractionToUintArray().0._State_11\, 
        \Unum::FractionToUintArray().0._State_12\);
    -- Signals:
    Signal \Unum::FractionToUintArray().0._Finished\: boolean := false;
    Signal \Unum::FractionToUintArray().0.return\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \Unum::FractionToUintArray().0.Unum::FractionWithHiddenBit().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::FractionToUintArray().0.Unum::FractionWithHiddenBit()._Started.0\: boolean := false;
    Signal \Unum::FractionToUintArray().0.Unum::ExponentValueWithBias().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::FractionToUintArray().0.Unum::ExponentValueWithBias()._Started.0\: boolean := false;
    Signal \Unum::FractionToUintArray().0.Unum::FractionSize().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::FractionToUintArray().0.Unum::FractionSize()._Started.0\: boolean := false;
    Signal \Unum::FractionToUintArray().0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::FractionToUintArray().0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Unum::FractionToUintArray().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\: boolean := false;
    Signal \Unum::FractionToUintArray().0.Unum::IsPositive().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::FractionToUintArray().0.Unum::IsPositive()._Started.0\: boolean := false;
    Signal \Unum::FractionToUintArray().0._Started\: boolean := false;
    Signal \Unum::FractionToUintArray().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::FractionToUintArray().0.Unum::FractionWithHiddenBit()._Finished.0\: boolean := false;
    Signal \Unum::FractionToUintArray().0.Unum::FractionWithHiddenBit().return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::FractionToUintArray().0.Unum::ExponentValueWithBias()._Finished.0\: boolean := false;
    Signal \Unum::FractionToUintArray().0.Unum::ExponentValueWithBias().return.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Unum::FractionToUintArray().0.Unum::FractionSize()._Finished.0\: boolean := false;
    Signal \Unum::FractionToUintArray().0.Unum::FractionSize().return.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::FractionToUintArray().0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\: boolean := false;
    Signal \Unum::FractionToUintArray().0.BitMask::op_LeftShift(BitMask,Int32).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::FractionToUintArray().0.Unum::IsPositive()._Finished.0\: boolean := false;
    Signal \Unum::FractionToUintArray().0.Unum::IsPositive().return.0\: boolean := false;
    -- System.UInt32[] Lombiq.Unum.Unum::FractionToUintArray().0 declarations end


    -- System.Boolean Lombiq.Unum.Unum::IsExact().0 declarations start
    -- State machine states:
    type \Unum::IsExact().0._States\ is (
        \Unum::IsExact().0._State_0\, 
        \Unum::IsExact().0._State_1\, 
        \Unum::IsExact().0._State_2\, 
        \Unum::IsExact().0._State_3\, 
        \Unum::IsExact().0._State_4\, 
        \Unum::IsExact().0._State_5\);
    -- Signals:
    Signal \Unum::IsExact().0._Finished\: boolean := false;
    Signal \Unum::IsExact().0.return\: boolean := false;
    Signal \Unum::IsExact().0.Unum::get_UncertaintyBitMask().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::IsExact().0.Unum::get_UncertaintyBitMask()._Started.0\: boolean := false;
    Signal \Unum::IsExact().0.BitMask::op_BitwiseAnd(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::IsExact().0.BitMask::op_BitwiseAnd(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::IsExact().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \Unum::IsExact().0.BitMask::op_Equality(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::IsExact().0.BitMask::op_Equality(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::IsExact().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \Unum::IsExact().0._Started\: boolean := false;
    Signal \Unum::IsExact().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::IsExact().0.Unum::get_UncertaintyBitMask()._Finished.0\: boolean := false;
    Signal \Unum::IsExact().0.Unum::get_UncertaintyBitMask().return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::IsExact().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \Unum::IsExact().0.BitMask::op_BitwiseAnd(BitMask,BitMask).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::IsExact().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \Unum::IsExact().0.BitMask::op_Equality(BitMask,BitMask).return.0\: boolean := false;
    -- System.Boolean Lombiq.Unum.Unum::IsExact().0 declarations end


    -- System.Boolean Lombiq.Unum.Unum::IsPositive().0 declarations start
    -- State machine states:
    type \Unum::IsPositive().0._States\ is (
        \Unum::IsPositive().0._State_0\, 
        \Unum::IsPositive().0._State_1\, 
        \Unum::IsPositive().0._State_2\, 
        \Unum::IsPositive().0._State_3\, 
        \Unum::IsPositive().0._State_4\, 
        \Unum::IsPositive().0._State_5\);
    -- Signals:
    Signal \Unum::IsPositive().0._Finished\: boolean := false;
    Signal \Unum::IsPositive().0.return\: boolean := false;
    Signal \Unum::IsPositive().0.Unum::get_SignBitMask().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::IsPositive().0.Unum::get_SignBitMask()._Started.0\: boolean := false;
    Signal \Unum::IsPositive().0.BitMask::op_BitwiseAnd(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::IsPositive().0.BitMask::op_BitwiseAnd(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::IsPositive().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \Unum::IsPositive().0.BitMask::op_Equality(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::IsPositive().0.BitMask::op_Equality(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::IsPositive().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \Unum::IsPositive().0._Started\: boolean := false;
    Signal \Unum::IsPositive().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::IsPositive().0.Unum::get_SignBitMask()._Finished.0\: boolean := false;
    Signal \Unum::IsPositive().0.Unum::get_SignBitMask().return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::IsPositive().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \Unum::IsPositive().0.BitMask::op_BitwiseAnd(BitMask,BitMask).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::IsPositive().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \Unum::IsPositive().0.BitMask::op_Equality(BitMask,BitMask).return.0\: boolean := false;
    -- System.Boolean Lombiq.Unum.Unum::IsPositive().0 declarations end


    -- System.Byte Lombiq.Unum.Unum::ExponentSize().0 declarations start
    -- State machine states:
    type \Unum::ExponentSize().0._States\ is (
        \Unum::ExponentSize().0._State_0\, 
        \Unum::ExponentSize().0._State_1\, 
        \Unum::ExponentSize().0._State_2\, 
        \Unum::ExponentSize().0._State_3\, 
        \Unum::ExponentSize().0._State_4\, 
        \Unum::ExponentSize().0._State_5\, 
        \Unum::ExponentSize().0._State_6\, 
        \Unum::ExponentSize().0._State_7\);
    -- Signals:
    Signal \Unum::ExponentSize().0._Finished\: boolean := false;
    Signal \Unum::ExponentSize().0.return\: unsigned(7 downto 0) := to_unsigned(0, 8);
    Signal \Unum::ExponentSize().0.Unum::get_ExponentSizeMask().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::ExponentSize().0.Unum::get_ExponentSizeMask()._Started.0\: boolean := false;
    Signal \Unum::ExponentSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \Unum::ExponentSize().0.BitMask::op_RightShift(BitMask,Int32).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentSize().0.BitMask::op_RightShift(BitMask,Int32).right.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Unum::ExponentSize().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\: boolean := false;
    Signal \Unum::ExponentSize().0.BitMask::op_Addition(BitMask,UInt32).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentSize().0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Unum::ExponentSize().0.BitMask::op_Addition(BitMask,UInt32)._Started.0\: boolean := false;
    Signal \Unum::ExponentSize().0.BitMask::GetLowest32Bits().this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentSize().0.BitMask::GetLowest32Bits()._Started.0\: boolean := false;
    Signal \Unum::ExponentSize().0._Started\: boolean := false;
    Signal \Unum::ExponentSize().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::ExponentSize().0.Unum::get_ExponentSizeMask()._Finished.0\: boolean := false;
    Signal \Unum::ExponentSize().0.Unum::get_ExponentSizeMask().return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \Unum::ExponentSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentSize().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\: boolean := false;
    Signal \Unum::ExponentSize().0.BitMask::op_RightShift(BitMask,Int32).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentSize().0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\: boolean := false;
    Signal \Unum::ExponentSize().0.BitMask::op_Addition(BitMask,UInt32).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentSize().0.BitMask::GetLowest32Bits()._Finished.0\: boolean := false;
    Signal \Unum::ExponentSize().0.BitMask::GetLowest32Bits().return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.Byte Lombiq.Unum.Unum::ExponentSize().0 declarations end


    -- System.UInt16 Lombiq.Unum.Unum::FractionSize().0 declarations start
    -- State machine states:
    type \Unum::FractionSize().0._States\ is (
        \Unum::FractionSize().0._State_0\, 
        \Unum::FractionSize().0._State_1\, 
        \Unum::FractionSize().0._State_2\, 
        \Unum::FractionSize().0._State_3\, 
        \Unum::FractionSize().0._State_4\, 
        \Unum::FractionSize().0._State_5\, 
        \Unum::FractionSize().0._State_6\);
    -- Signals:
    Signal \Unum::FractionSize().0._Finished\: boolean := false;
    Signal \Unum::FractionSize().0.return\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::FractionSize().0.Unum::get_FractionSizeMask().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::FractionSize().0.Unum::get_FractionSizeMask()._Started.0\: boolean := false;
    Signal \Unum::FractionSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::FractionSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::FractionSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \Unum::FractionSize().0.BitMask::op_Addition(BitMask,UInt32).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::FractionSize().0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Unum::FractionSize().0.BitMask::op_Addition(BitMask,UInt32)._Started.0\: boolean := false;
    Signal \Unum::FractionSize().0.BitMask::GetLowest32Bits().this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::FractionSize().0.BitMask::GetLowest32Bits()._Started.0\: boolean := false;
    Signal \Unum::FractionSize().0._Started\: boolean := false;
    Signal \Unum::FractionSize().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::FractionSize().0.Unum::get_FractionSizeMask()._Finished.0\: boolean := false;
    Signal \Unum::FractionSize().0.Unum::get_FractionSizeMask().return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::FractionSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \Unum::FractionSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::FractionSize().0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\: boolean := false;
    Signal \Unum::FractionSize().0.BitMask::op_Addition(BitMask,UInt32).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::FractionSize().0.BitMask::GetLowest32Bits()._Finished.0\: boolean := false;
    Signal \Unum::FractionSize().0.BitMask::GetLowest32Bits().return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.UInt16 Lombiq.Unum.Unum::FractionSize().0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionMask().0 declarations start
    -- State machine states:
    type \Unum::FractionMask().0._States\ is (
        \Unum::FractionMask().0._State_0\, 
        \Unum::FractionMask().0._State_1\, 
        \Unum::FractionMask().0._State_2\, 
        \Unum::FractionMask().0._State_3\, 
        \Unum::FractionMask().0._State_4\, 
        \Unum::FractionMask().0._State_5\, 
        \Unum::FractionMask().0._State_6\, 
        \Unum::FractionMask().0._State_7\, 
        \Unum::FractionMask().0._State_8\, 
        \Unum::FractionMask().0._State_9\);
    -- Signals:
    Signal \Unum::FractionMask().0._Finished\: boolean := false;
    Signal \Unum::FractionMask().0.return\: \Lombiq.Unum.BitMask\;
    Signal \Unum::FractionMask().0.Unum::get_Size().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::FractionMask().0.Unum::get_Size()._Started.0\: boolean := false;
    Signal \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16)._Started.0\: boolean := false;
    Signal \Unum::FractionMask().0.Unum::FractionSize()._Started.0\: boolean := false;
    Signal \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\: boolean := false;
    Signal \Unum::FractionMask().0.BitMask::op_Subtraction(BitMask,UInt32).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::FractionMask().0.BitMask::op_Subtraction(BitMask,UInt32).right.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Unum::FractionMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\: boolean := false;
    Signal \Unum::FractionMask().0._Started\: boolean := false;
    Signal \Unum::FractionMask().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::FractionMask().0.Unum::get_Size()._Finished.0\: boolean := false;
    Signal \Unum::FractionMask().0.Unum::get_Size().return.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\: boolean := false;
    Signal \Unum::FractionMask().0.Unum::FractionSize()._Finished.0\: boolean := false;
    Signal \Unum::FractionMask().0.Unum::FractionSize().return.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\: boolean := false;
    Signal \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::FractionMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\: boolean := false;
    Signal \Unum::FractionMask().0.BitMask::op_Subtraction(BitMask,UInt32).return.0\: \Lombiq.Unum.BitMask\;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionMask().0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentMask().0 declarations start
    -- State machine states:
    type \Unum::ExponentMask().0._States\ is (
        \Unum::ExponentMask().0._State_0\, 
        \Unum::ExponentMask().0._State_1\, 
        \Unum::ExponentMask().0._State_2\, 
        \Unum::ExponentMask().0._State_3\, 
        \Unum::ExponentMask().0._State_4\, 
        \Unum::ExponentMask().0._State_5\, 
        \Unum::ExponentMask().0._State_6\, 
        \Unum::ExponentMask().0._State_7\, 
        \Unum::ExponentMask().0._State_8\, 
        \Unum::ExponentMask().0._State_9\);
    -- Signals:
    Signal \Unum::ExponentMask().0._Finished\: boolean := false;
    Signal \Unum::ExponentMask().0.return\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentMask().0.Unum::get_Size().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::ExponentMask().0.Unum::get_Size()._Started.0\: boolean := false;
    Signal \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16)._Started.0\: boolean := false;
    Signal \Unum::ExponentMask().0.Unum::ExponentSize()._Started.0\: boolean := false;
    Signal \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\: boolean := false;
    Signal \Unum::ExponentMask().0.BitMask::op_Subtraction(BitMask,UInt32).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentMask().0.BitMask::op_Subtraction(BitMask,UInt32).right.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Unum::ExponentMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\: boolean := false;
    Signal \Unum::ExponentMask().0.Unum::FractionSize()._Started.0\: boolean := false;
    Signal \Unum::ExponentMask().0._Started\: boolean := false;
    Signal \Unum::ExponentMask().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::ExponentMask().0.Unum::get_Size()._Finished.0\: boolean := false;
    Signal \Unum::ExponentMask().0.Unum::get_Size().return.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\: boolean := false;
    Signal \Unum::ExponentMask().0.Unum::ExponentSize()._Finished.0\: boolean := false;
    Signal \Unum::ExponentMask().0.Unum::ExponentSize().return.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
    Signal \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\: boolean := false;
    Signal \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\: boolean := false;
    Signal \Unum::ExponentMask().0.BitMask::op_Subtraction(BitMask,UInt32).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentMask().0.Unum::FractionSize()._Finished.0\: boolean := false;
    Signal \Unum::ExponentMask().0.Unum::FractionSize().return.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentMask().0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::Exponent().0 declarations start
    -- State machine states:
    type \Unum::Exponent().0._States\ is (
        \Unum::Exponent().0._State_0\, 
        \Unum::Exponent().0._State_1\, 
        \Unum::Exponent().0._State_2\, 
        \Unum::Exponent().0._State_3\, 
        \Unum::Exponent().0._State_4\, 
        \Unum::Exponent().0._State_5\, 
        \Unum::Exponent().0._State_6\);
    -- Signals:
    Signal \Unum::Exponent().0._Finished\: boolean := false;
    Signal \Unum::Exponent().0.return\: \Lombiq.Unum.BitMask\;
    Signal \Unum::Exponent().0.Unum::ExponentMask()._Started.0\: boolean := false;
    Signal \Unum::Exponent().0.BitMask::op_BitwiseAnd(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::Exponent().0.BitMask::op_BitwiseAnd(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::Exponent().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \Unum::Exponent().0.Unum::FractionSize()._Started.0\: boolean := false;
    Signal \Unum::Exponent().0.BitMask::op_RightShift(BitMask,Int32).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::Exponent().0.BitMask::op_RightShift(BitMask,Int32).right.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Unum::Exponent().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\: boolean := false;
    Signal \Unum::Exponent().0._Started\: boolean := false;
    Signal \Unum::Exponent().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::Exponent().0.Unum::ExponentMask()._Finished.0\: boolean := false;
    Signal \Unum::Exponent().0.Unum::ExponentMask().return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::Exponent().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \Unum::Exponent().0.BitMask::op_BitwiseAnd(BitMask,BitMask).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::Exponent().0.Unum::FractionSize()._Finished.0\: boolean := false;
    Signal \Unum::Exponent().0.Unum::FractionSize().return.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::Exponent().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\: boolean := false;
    Signal \Unum::Exponent().0.BitMask::op_RightShift(BitMask,Int32).return.0\: \Lombiq.Unum.BitMask\;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::Exponent().0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::Fraction().0 declarations start
    -- State machine states:
    type \Unum::Fraction().0._States\ is (
        \Unum::Fraction().0._State_0\, 
        \Unum::Fraction().0._State_1\, 
        \Unum::Fraction().0._State_2\, 
        \Unum::Fraction().0._State_3\, 
        \Unum::Fraction().0._State_4\, 
        \Unum::Fraction().0._State_5\);
    -- Signals:
    Signal \Unum::Fraction().0._Finished\: boolean := false;
    Signal \Unum::Fraction().0.return\: \Lombiq.Unum.BitMask\;
    Signal \Unum::Fraction().0.Unum::FractionMask()._Started.0\: boolean := false;
    Signal \Unum::Fraction().0.BitMask::op_BitwiseAnd(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::Fraction().0.BitMask::op_BitwiseAnd(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::Fraction().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \Unum::Fraction().0.BitMask::op_RightShift(BitMask,Int32).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::Fraction().0.BitMask::op_RightShift(BitMask,Int32).right.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Unum::Fraction().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\: boolean := false;
    Signal \Unum::Fraction().0._Started\: boolean := false;
    Signal \Unum::Fraction().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::Fraction().0.Unum::FractionMask()._Finished.0\: boolean := false;
    Signal \Unum::Fraction().0.Unum::FractionMask().return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::Fraction().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \Unum::Fraction().0.BitMask::op_BitwiseAnd(BitMask,BitMask).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::Fraction().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\: boolean := false;
    Signal \Unum::Fraction().0.BitMask::op_RightShift(BitMask,Int32).return.0\: \Lombiq.Unum.BitMask\;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::Fraction().0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit().0 declarations start
    -- State machine states:
    type \Unum::FractionWithHiddenBit().0._States\ is (
        \Unum::FractionWithHiddenBit().0._State_0\, 
        \Unum::FractionWithHiddenBit().0._State_1\, 
        \Unum::FractionWithHiddenBit().0._State_2\, 
        \Unum::FractionWithHiddenBit().0._State_3\, 
        \Unum::FractionWithHiddenBit().0._State_4\, 
        \Unum::FractionWithHiddenBit().0._State_5\, 
        \Unum::FractionWithHiddenBit().0._State_6\, 
        \Unum::FractionWithHiddenBit().0._State_7\, 
        \Unum::FractionWithHiddenBit().0._State_8\, 
        \Unum::FractionWithHiddenBit().0._State_9\, 
        \Unum::FractionWithHiddenBit().0._State_10\);
    -- Signals:
    Signal \Unum::FractionWithHiddenBit().0._Finished\: boolean := false;
    Signal \Unum::FractionWithHiddenBit().0.return\: \Lombiq.Unum.BitMask\;
    Signal \Unum::FractionWithHiddenBit().0.Unum::HiddenBitIsOne().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::FractionWithHiddenBit().0.Unum::HiddenBitIsOne()._Started.0\: boolean := false;
    Signal \Unum::FractionWithHiddenBit().0.Unum::Fraction()._Started.0\: boolean := false;
    Signal \Unum::FractionWithHiddenBit().0.Unum::FractionSize()._Started.0\: boolean := false;
    Signal \Unum::FractionWithHiddenBit().0.BitMask::SetOne(UInt16).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::FractionWithHiddenBit().0.BitMask::SetOne(UInt16).index.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::FractionWithHiddenBit().0.BitMask::SetOne(UInt16)._Started.0\: boolean := false;
    Signal \Unum::FractionWithHiddenBit().0._Started\: boolean := false;
    Signal \Unum::FractionWithHiddenBit().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::FractionWithHiddenBit().0.Unum::HiddenBitIsOne()._Finished.0\: boolean := false;
    Signal \Unum::FractionWithHiddenBit().0.Unum::HiddenBitIsOne().return.0\: boolean := false;
    Signal \Unum::FractionWithHiddenBit().0.Unum::Fraction()._Finished.0\: boolean := false;
    Signal \Unum::FractionWithHiddenBit().0.Unum::Fraction().return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::FractionWithHiddenBit().0.Unum::FractionSize()._Finished.0\: boolean := false;
    Signal \Unum::FractionWithHiddenBit().0.Unum::FractionSize().return.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::FractionWithHiddenBit().0.BitMask::SetOne(UInt16)._Finished.0\: boolean := false;
    Signal \Unum::FractionWithHiddenBit().0.BitMask::SetOne(UInt16).return.0\: \Lombiq.Unum.BitMask\;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit().0 declarations end


    -- System.Int32 Lombiq.Unum.Unum::Bias().0 declarations start
    -- State machine states:
    type \Unum::Bias().0._States\ is (
        \Unum::Bias().0._State_0\, 
        \Unum::Bias().0._State_1\, 
        \Unum::Bias().0._State_2\, 
        \Unum::Bias().0._State_3\);
    -- Signals:
    Signal \Unum::Bias().0._Finished\: boolean := false;
    Signal \Unum::Bias().0.return\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Unum::Bias().0.Unum::ExponentSize()._Started.0\: boolean := false;
    Signal \Unum::Bias().0._Started\: boolean := false;
    Signal \Unum::Bias().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::Bias().0.Unum::ExponentSize()._Finished.0\: boolean := false;
    Signal \Unum::Bias().0.Unum::ExponentSize().return.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
    -- System.Int32 Lombiq.Unum.Unum::Bias().0 declarations end


    -- System.Boolean Lombiq.Unum.Unum::HiddenBitIsOne().0 declarations start
    -- State machine states:
    type \Unum::HiddenBitIsOne().0._States\ is (
        \Unum::HiddenBitIsOne().0._State_0\, 
        \Unum::HiddenBitIsOne().0._State_1\, 
        \Unum::HiddenBitIsOne().0._State_2\, 
        \Unum::HiddenBitIsOne().0._State_3\, 
        \Unum::HiddenBitIsOne().0._State_4\);
    -- Signals:
    Signal \Unum::HiddenBitIsOne().0._Finished\: boolean := false;
    Signal \Unum::HiddenBitIsOne().0.return\: boolean := false;
    Signal \Unum::HiddenBitIsOne().0.Unum::Exponent()._Started.0\: boolean := false;
    Signal \Unum::HiddenBitIsOne().0.BitMask::GetLowest32Bits().this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::HiddenBitIsOne().0.BitMask::GetLowest32Bits()._Started.0\: boolean := false;
    Signal \Unum::HiddenBitIsOne().0._Started\: boolean := false;
    Signal \Unum::HiddenBitIsOne().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::HiddenBitIsOne().0.Unum::Exponent()._Finished.0\: boolean := false;
    Signal \Unum::HiddenBitIsOne().0.Unum::Exponent().return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::HiddenBitIsOne().0.BitMask::GetLowest32Bits()._Finished.0\: boolean := false;
    Signal \Unum::HiddenBitIsOne().0.BitMask::GetLowest32Bits().return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.Boolean Lombiq.Unum.Unum::HiddenBitIsOne().0 declarations end


    -- System.Int32 Lombiq.Unum.Unum::ExponentValueWithBias().0 declarations start
    -- State machine states:
    type \Unum::ExponentValueWithBias().0._States\ is (
        \Unum::ExponentValueWithBias().0._State_0\, 
        \Unum::ExponentValueWithBias().0._State_1\, 
        \Unum::ExponentValueWithBias().0._State_2\, 
        \Unum::ExponentValueWithBias().0._State_3\, 
        \Unum::ExponentValueWithBias().0._State_4\, 
        \Unum::ExponentValueWithBias().0._State_5\, 
        \Unum::ExponentValueWithBias().0._State_6\, 
        \Unum::ExponentValueWithBias().0._State_7\, 
        \Unum::ExponentValueWithBias().0._State_8\, 
        \Unum::ExponentValueWithBias().0._State_9\);
    -- Signals:
    Signal \Unum::ExponentValueWithBias().0._Finished\: boolean := false;
    Signal \Unum::ExponentValueWithBias().0.return\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Unum::ExponentValueWithBias().0.Unum::HiddenBitIsOne()._Started.0\: boolean := false;
    Signal \Unum::ExponentValueWithBias().0.Unum::Exponent()._Started.0\: boolean := false;
    Signal \Unum::ExponentValueWithBias().0.BitMask::GetLowest32Bits().this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentValueWithBias().0.BitMask::GetLowest32Bits()._Started.0\: boolean := false;
    Signal \Unum::ExponentValueWithBias().0.Unum::Bias()._Started.0\: boolean := false;
    Signal \Unum::ExponentValueWithBias().0._Started\: boolean := false;
    Signal \Unum::ExponentValueWithBias().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::ExponentValueWithBias().0.Unum::HiddenBitIsOne()._Finished.0\: boolean := false;
    Signal \Unum::ExponentValueWithBias().0.Unum::HiddenBitIsOne().return.0\: boolean := false;
    Signal \Unum::ExponentValueWithBias().0.Unum::Exponent()._Finished.0\: boolean := false;
    Signal \Unum::ExponentValueWithBias().0.Unum::Exponent().return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentValueWithBias().0.BitMask::GetLowest32Bits()._Finished.0\: boolean := false;
    Signal \Unum::ExponentValueWithBias().0.BitMask::GetLowest32Bits().return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Unum::ExponentValueWithBias().0.Unum::Bias()._Finished.0\: boolean := false;
    Signal \Unum::ExponentValueWithBias().0.Unum::Bias().return.0\: signed(31 downto 0) := to_signed(0, 32);
    -- System.Int32 Lombiq.Unum.Unum::ExponentValueWithBias().0 declarations end


    -- System.Boolean Lombiq.Unum.Unum::IsNan().0 declarations start
    -- State machine states:
    type \Unum::IsNan().0._States\ is (
        \Unum::IsNan().0._State_0\, 
        \Unum::IsNan().0._State_1\, 
        \Unum::IsNan().0._State_2\, 
        \Unum::IsNan().0._State_3\, 
        \Unum::IsNan().0._State_4\, 
        \Unum::IsNan().0._State_5\, 
        \Unum::IsNan().0._State_6\, 
        \Unum::IsNan().0._State_7\);
    -- Signals:
    Signal \Unum::IsNan().0._Finished\: boolean := false;
    Signal \Unum::IsNan().0.return\: boolean := false;
    Signal \Unum::IsNan().0.Unum::get_SignalingNotANumber().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::IsNan().0.Unum::get_SignalingNotANumber()._Started.0\: boolean := false;
    Signal \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \Unum::IsNan().0.Unum::get_QuietNotANumber().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::IsNan().0.Unum::get_QuietNotANumber()._Started.0\: boolean := false;
    Signal \Unum::IsNan().0._Started\: boolean := false;
    Signal \Unum::IsNan().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::IsNan().0.Unum::get_SignalingNotANumber()._Finished.0\: boolean := false;
    Signal \Unum::IsNan().0.Unum::get_SignalingNotANumber().return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask).return.0\: boolean := false;
    Signal \Unum::IsNan().0.Unum::get_QuietNotANumber()._Finished.0\: boolean := false;
    Signal \Unum::IsNan().0.Unum::get_QuietNotANumber().return.0\: \Lombiq.Unum.BitMask\;
    -- System.Boolean Lombiq.Unum.Unum::IsNan().0 declarations end


    -- System.Boolean Lombiq.Unum.Unum::IsPositiveInfinity().0 declarations start
    -- State machine states:
    type \Unum::IsPositiveInfinity().0._States\ is (
        \Unum::IsPositiveInfinity().0._State_0\, 
        \Unum::IsPositiveInfinity().0._State_1\, 
        \Unum::IsPositiveInfinity().0._State_2\, 
        \Unum::IsPositiveInfinity().0._State_3\, 
        \Unum::IsPositiveInfinity().0._State_4\);
    -- Signals:
    Signal \Unum::IsPositiveInfinity().0._Finished\: boolean := false;
    Signal \Unum::IsPositiveInfinity().0.return\: boolean := false;
    Signal \Unum::IsPositiveInfinity().0.Unum::get_PositiveInfinity().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::IsPositiveInfinity().0.Unum::get_PositiveInfinity()._Started.0\: boolean := false;
    Signal \Unum::IsPositiveInfinity().0.BitMask::op_Equality(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::IsPositiveInfinity().0.BitMask::op_Equality(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::IsPositiveInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \Unum::IsPositiveInfinity().0._Started\: boolean := false;
    Signal \Unum::IsPositiveInfinity().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::IsPositiveInfinity().0.Unum::get_PositiveInfinity()._Finished.0\: boolean := false;
    Signal \Unum::IsPositiveInfinity().0.Unum::get_PositiveInfinity().return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::IsPositiveInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \Unum::IsPositiveInfinity().0.BitMask::op_Equality(BitMask,BitMask).return.0\: boolean := false;
    -- System.Boolean Lombiq.Unum.Unum::IsPositiveInfinity().0 declarations end


    -- System.Boolean Lombiq.Unum.Unum::IsNegativeInfinity().0 declarations start
    -- State machine states:
    type \Unum::IsNegativeInfinity().0._States\ is (
        \Unum::IsNegativeInfinity().0._State_0\, 
        \Unum::IsNegativeInfinity().0._State_1\, 
        \Unum::IsNegativeInfinity().0._State_2\, 
        \Unum::IsNegativeInfinity().0._State_3\, 
        \Unum::IsNegativeInfinity().0._State_4\);
    -- Signals:
    Signal \Unum::IsNegativeInfinity().0._Finished\: boolean := false;
    Signal \Unum::IsNegativeInfinity().0.return\: boolean := false;
    Signal \Unum::IsNegativeInfinity().0.Unum::get_NegativeInfinity().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::IsNegativeInfinity().0.Unum::get_NegativeInfinity()._Started.0\: boolean := false;
    Signal \Unum::IsNegativeInfinity().0.BitMask::op_Equality(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::IsNegativeInfinity().0.BitMask::op_Equality(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::IsNegativeInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \Unum::IsNegativeInfinity().0._Started\: boolean := false;
    Signal \Unum::IsNegativeInfinity().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::IsNegativeInfinity().0.Unum::get_NegativeInfinity()._Finished.0\: boolean := false;
    Signal \Unum::IsNegativeInfinity().0.Unum::get_NegativeInfinity().return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::IsNegativeInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \Unum::IsNegativeInfinity().0.BitMask::op_Equality(BitMask,BitMask).return.0\: boolean := false;
    -- System.Boolean Lombiq.Unum.Unum::IsNegativeInfinity().0 declarations end


    -- Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0 declarations start
    -- State machine states:
    type \Unum::AddExactUnums(Unum,Unum).0._States\ is (
        \Unum::AddExactUnums(Unum,Unum).0._State_0\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_1\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_2\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_3\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_4\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_5\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_6\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_7\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_8\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_9\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_10\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_11\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_12\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_13\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_14\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_15\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_16\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_17\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_18\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_19\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_20\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_21\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_22\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_23\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_24\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_25\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_26\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_27\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_28\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_29\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_30\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_31\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_32\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_33\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_34\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_35\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_36\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_37\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_38\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_39\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_40\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_41\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_42\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_43\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_44\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_45\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_46\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_47\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_48\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_49\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_50\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_51\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_52\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_53\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_54\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_55\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_56\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_57\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_58\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_59\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_60\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_61\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_62\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_63\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_64\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_65\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_66\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_67\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_68\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_69\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_70\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_71\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_72\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_73\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_74\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_75\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_76\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_77\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_78\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_79\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_80\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_81\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_82\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_83\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_84\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_85\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_86\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_87\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_88\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_89\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_90\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_91\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_92\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_93\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_94\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_95\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_96\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_97\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_98\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_99\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_100\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_101\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_102\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_103\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_104\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_105\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_106\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_107\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_108\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_109\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_110\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_111\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_112\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_113\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_114\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_115\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_116\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_117\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_118\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_119\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_120\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_121\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_122\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_123\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_124\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_125\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_126\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_127\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_128\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_129\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_130\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_131\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_132\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_133\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_134\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_135\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_136\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_137\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_138\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_139\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_140\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_141\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_142\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_143\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_144\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_145\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_146\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_147\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_148\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_149\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_150\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_151\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_152\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_153\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_154\, 
        \Unum::AddExactUnums(Unum,Unum).0._State_155\);
    -- Signals:
    Signal \Unum::AddExactUnums(Unum,Unum).0._Finished\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.return\: \Lombiq.Unum.Unum\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean)._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNan().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNan()._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber()._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).environment.parameter.Out.0\: \Lombiq.Unum.UnumEnvironment\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).bits.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask)._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity()._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity()._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::get_PositiveInfinity().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::get_PositiveInfinity()._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::get_NegativeInfinity().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::get_NegativeInfinity()._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment).this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment).environment.parameter.Out.0\: \Lombiq.Unum.UnumEnvironment\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment)._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean).signBitsMatch.parameter.Out.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean)._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne()._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction()._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_GreaterThanOrEqual(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_GreaterThanOrEqual(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_GreaterThanOrEqual(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition().this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::get_Size().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::get_Size()._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueToExponentBits(Int32,Byte).value.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueToExponentBits(Int32,Byte).size.parameter.Out.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueToExponentBits(Int32,Byte)._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_Addition(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_Addition(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::ShiftOutLeastSignificantZeros().this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::ShiftOutLeastSignificantZeros()._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::SetZero(UInt16).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::SetZero(UInt16).index.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::SetZero(UInt16)._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::IsExact().this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::IsExact()._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).this.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).signBit.parameter.Out.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).exponent.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).fraction.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).uncertainityBit.parameter.Out.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).exponentSize.parameter.Out.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).fractionSize.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Started.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0._Started\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.left.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.right.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNan()._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNan().return.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber()._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber().return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).this.parameter.In.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).environment.parameter.In.0\: \Lombiq.Unum.UnumEnvironment\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask)._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity()._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity().return.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity()._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity().return.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::get_PositiveInfinity()._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::get_PositiveInfinity().return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::get_NegativeInfinity()._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::get_NegativeInfinity().return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment).this.parameter.In.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment).environment.parameter.In.0\: \Lombiq.Unum.UnumEnvironment\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment)._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias().return.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive().return.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax().return.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize().return.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit().return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean)._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne()._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne().return.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction()._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction().return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_GreaterThanOrEqual(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_GreaterThanOrEqual(BitMask,BitMask).return.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition().return.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::get_Size()._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::get_Size().return.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueToExponentBits(Int32,Byte)._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueToExponentBits(Int32,Byte).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_Addition(BitMask,BitMask).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::ShiftOutLeastSignificantZeros()._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::ShiftOutLeastSignificantZeros().return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::SetZero(UInt16)._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.BitMask::SetZero(UInt16).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::IsExact()._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::IsExact().return.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Finished.0\: boolean := false;
    Signal \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).return.0\: \Lombiq.Unum.BitMask\;
    -- Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentValueToExponentBits(System.Int32,System.Byte).0 declarations start
    -- State machine states:
    type \Unum::ExponentValueToExponentBits(Int32,Byte).0._States\ is (
        \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_0\, 
        \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_1\, 
        \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_2\, 
        \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_3\, 
        \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_4\, 
        \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_5\, 
        \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_6\, 
        \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_7\, 
        \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_8\, 
        \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_9\, 
        \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_10\);
    -- Signals:
    Signal \Unum::ExponentValueToExponentBits(Int32,Byte).0._Finished\: boolean := false;
    Signal \Unum::ExponentValueToExponentBits(Int32,Byte).0.return\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\: boolean := false;
    Signal \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\: boolean := false;
    Signal \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).right.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\: boolean := false;
    Signal \Unum::ExponentValueToExponentBits(Int32,Byte).0._Started\: boolean := false;
    Signal \Unum::ExponentValueToExponentBits(Int32,Byte).0.value.parameter.In\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Unum::ExponentValueToExponentBits(Int32,Byte).0.size.parameter.In\: unsigned(7 downto 0) := to_unsigned(0, 8);
    Signal \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
    Signal \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\: boolean := false;
    Signal \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\: boolean := false;
    Signal \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\: boolean := false;
    Signal \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).return.0\: \Lombiq.Unum.BitMask\;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentValueToExponentBits(System.Int32,System.Byte).0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::AddAlignedFractions(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean).0 declarations start
    -- State machine states:
    type \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._States\ is (
        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_0\, 
        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_1\, 
        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_2\, 
        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_3\, 
        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_4\, 
        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_5\, 
        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_6\, 
        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_7\, 
        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_8\, 
        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_9\, 
        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_10\, 
        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_11\, 
        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_12\, 
        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_13\, 
        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_14\);
    -- Signals:
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._Finished\: boolean := false;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.return\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\: boolean := false;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean)._Started.0\: boolean := false;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Addition(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Addition(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_GreaterThan(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_GreaterThan(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_GreaterThan(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._Started\: boolean := false;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.left.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.right.parameter.In\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.signBitsMatch.parameter.In\: boolean := false;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\: boolean := false;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Addition(BitMask,BitMask).return.0\: \Lombiq.Unum.BitMask\;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_GreaterThan(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_GreaterThan(BitMask,BitMask).return.0\: boolean := false;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask).return.0\: \Lombiq.Unum.BitMask\;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::AddAlignedFractions(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean).0 declarations end


    -- Lombiq.Unum.Unum Lombiq.Unum.Unum::op_Addition(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0 declarations start
    -- State machine states:
    type \Unum::op_Addition(Unum,Unum).0._States\ is (
        \Unum::op_Addition(Unum,Unum).0._State_0\, 
        \Unum::op_Addition(Unum,Unum).0._State_1\, 
        \Unum::op_Addition(Unum,Unum).0._State_2\, 
        \Unum::op_Addition(Unum,Unum).0._State_3\);
    -- Signals:
    Signal \Unum::op_Addition(Unum,Unum).0._Finished\: boolean := false;
    Signal \Unum::op_Addition(Unum,Unum).0.return\: \Lombiq.Unum.Unum\;
    Signal \Unum::op_Addition(Unum,Unum).0.Unum::AddExactUnums(Unum,Unum).left.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::op_Addition(Unum,Unum).0.Unum::AddExactUnums(Unum,Unum).right.parameter.Out.0\: \Lombiq.Unum.Unum\;
    Signal \Unum::op_Addition(Unum,Unum).0.Unum::AddExactUnums(Unum,Unum)._Started.0\: boolean := false;
    Signal \Unum::op_Addition(Unum,Unum).0._Started\: boolean := false;
    Signal \Unum::op_Addition(Unum,Unum).0.left.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::op_Addition(Unum,Unum).0.right.parameter.In\: \Lombiq.Unum.Unum\;
    Signal \Unum::op_Addition(Unum,Unum).0.Unum::AddExactUnums(Unum,Unum)._Finished.0\: boolean := false;
    Signal \Unum::op_Addition(Unum,Unum).0.Unum::AddExactUnums(Unum,Unum).return.0\: \Lombiq.Unum.Unum\;
    -- Lombiq.Unum.Unum Lombiq.Unum.Unum::op_Addition(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0 declarations end


    -- System.UInt16 Lombiq.Unum.Unum::get_FractionSizeMax().0 declarations start
    -- State machine states:
    type \Unum::get_FractionSizeMax().0._States\ is (
        \Unum::get_FractionSizeMax().0._State_0\, 
        \Unum::get_FractionSizeMax().0._State_1\, 
        \Unum::get_FractionSizeMax().0._State_2\);
    -- Signals:
    Signal \Unum::get_FractionSizeMax().0._Finished\: boolean := false;
    Signal \Unum::get_FractionSizeMax().0.return\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::get_FractionSizeMax().0._Started\: boolean := false;
    Signal \Unum::get_FractionSizeMax().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    -- System.UInt16 Lombiq.Unum.Unum::get_FractionSizeMax().0 declarations end


    -- System.UInt16 Lombiq.Unum.Unum::get_Size().0 declarations start
    -- State machine states:
    type \Unum::get_Size().0._States\ is (
        \Unum::get_Size().0._State_0\, 
        \Unum::get_Size().0._State_1\, 
        \Unum::get_Size().0._State_2\);
    -- Signals:
    Signal \Unum::get_Size().0._Finished\: boolean := false;
    Signal \Unum::get_Size().0.return\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Unum::get_Size().0._Started\: boolean := false;
    Signal \Unum::get_Size().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    -- System.UInt16 Lombiq.Unum.Unum::get_Size().0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_UncertaintyBitMask().0 declarations start
    -- State machine states:
    type \Unum::get_UncertaintyBitMask().0._States\ is (
        \Unum::get_UncertaintyBitMask().0._State_0\, 
        \Unum::get_UncertaintyBitMask().0._State_1\, 
        \Unum::get_UncertaintyBitMask().0._State_2\);
    -- Signals:
    Signal \Unum::get_UncertaintyBitMask().0._Finished\: boolean := false;
    Signal \Unum::get_UncertaintyBitMask().0.return\: \Lombiq.Unum.BitMask\;
    Signal \Unum::get_UncertaintyBitMask().0._Started\: boolean := false;
    Signal \Unum::get_UncertaintyBitMask().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_UncertaintyBitMask().0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_ExponentSizeMask().0 declarations start
    -- State machine states:
    type \Unum::get_ExponentSizeMask().0._States\ is (
        \Unum::get_ExponentSizeMask().0._State_0\, 
        \Unum::get_ExponentSizeMask().0._State_1\, 
        \Unum::get_ExponentSizeMask().0._State_2\);
    -- Signals:
    Signal \Unum::get_ExponentSizeMask().0._Finished\: boolean := false;
    Signal \Unum::get_ExponentSizeMask().0.return\: \Lombiq.Unum.BitMask\;
    Signal \Unum::get_ExponentSizeMask().0._Started\: boolean := false;
    Signal \Unum::get_ExponentSizeMask().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_ExponentSizeMask().0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_FractionSizeMask().0 declarations start
    -- State machine states:
    type \Unum::get_FractionSizeMask().0._States\ is (
        \Unum::get_FractionSizeMask().0._State_0\, 
        \Unum::get_FractionSizeMask().0._State_1\, 
        \Unum::get_FractionSizeMask().0._State_2\);
    -- Signals:
    Signal \Unum::get_FractionSizeMask().0._Finished\: boolean := false;
    Signal \Unum::get_FractionSizeMask().0.return\: \Lombiq.Unum.BitMask\;
    Signal \Unum::get_FractionSizeMask().0._Started\: boolean := false;
    Signal \Unum::get_FractionSizeMask().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_FractionSizeMask().0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_SignBitMask().0 declarations start
    -- State machine states:
    type \Unum::get_SignBitMask().0._States\ is (
        \Unum::get_SignBitMask().0._State_0\, 
        \Unum::get_SignBitMask().0._State_1\, 
        \Unum::get_SignBitMask().0._State_2\);
    -- Signals:
    Signal \Unum::get_SignBitMask().0._Finished\: boolean := false;
    Signal \Unum::get_SignBitMask().0.return\: \Lombiq.Unum.BitMask\;
    Signal \Unum::get_SignBitMask().0._Started\: boolean := false;
    Signal \Unum::get_SignBitMask().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_SignBitMask().0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_PositiveInfinity().0 declarations start
    -- State machine states:
    type \Unum::get_PositiveInfinity().0._States\ is (
        \Unum::get_PositiveInfinity().0._State_0\, 
        \Unum::get_PositiveInfinity().0._State_1\, 
        \Unum::get_PositiveInfinity().0._State_2\);
    -- Signals:
    Signal \Unum::get_PositiveInfinity().0._Finished\: boolean := false;
    Signal \Unum::get_PositiveInfinity().0.return\: \Lombiq.Unum.BitMask\;
    Signal \Unum::get_PositiveInfinity().0._Started\: boolean := false;
    Signal \Unum::get_PositiveInfinity().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_PositiveInfinity().0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_NegativeInfinity().0 declarations start
    -- State machine states:
    type \Unum::get_NegativeInfinity().0._States\ is (
        \Unum::get_NegativeInfinity().0._State_0\, 
        \Unum::get_NegativeInfinity().0._State_1\, 
        \Unum::get_NegativeInfinity().0._State_2\);
    -- Signals:
    Signal \Unum::get_NegativeInfinity().0._Finished\: boolean := false;
    Signal \Unum::get_NegativeInfinity().0.return\: \Lombiq.Unum.BitMask\;
    Signal \Unum::get_NegativeInfinity().0._Started\: boolean := false;
    Signal \Unum::get_NegativeInfinity().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_NegativeInfinity().0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_QuietNotANumber().0 declarations start
    -- State machine states:
    type \Unum::get_QuietNotANumber().0._States\ is (
        \Unum::get_QuietNotANumber().0._State_0\, 
        \Unum::get_QuietNotANumber().0._State_1\, 
        \Unum::get_QuietNotANumber().0._State_2\);
    -- Signals:
    Signal \Unum::get_QuietNotANumber().0._Finished\: boolean := false;
    Signal \Unum::get_QuietNotANumber().0.return\: \Lombiq.Unum.BitMask\;
    Signal \Unum::get_QuietNotANumber().0._Started\: boolean := false;
    Signal \Unum::get_QuietNotANumber().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_QuietNotANumber().0 declarations end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_SignalingNotANumber().0 declarations start
    -- State machine states:
    type \Unum::get_SignalingNotANumber().0._States\ is (
        \Unum::get_SignalingNotANumber().0._State_0\, 
        \Unum::get_SignalingNotANumber().0._State_1\, 
        \Unum::get_SignalingNotANumber().0._State_2\);
    -- Signals:
    Signal \Unum::get_SignalingNotANumber().0._Finished\: boolean := false;
    Signal \Unum::get_SignalingNotANumber().0.return\: \Lombiq.Unum.BitMask\;
    Signal \Unum::get_SignalingNotANumber().0._Started\: boolean := false;
    Signal \Unum::get_SignalingNotANumber().0.this.parameter.In\: \Lombiq.Unum.Unum\;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_SignalingNotANumber().0 declarations end


    -- System.UInt16 Lombiq.Unum.UnumHelper::SegmentSizeSizeToSegmentSize(System.Byte).0 declarations start
    -- State machine states:
    type \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._States\ is (
        \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._State_0\, 
        \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._State_1\, 
        \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._State_2\);
    -- Signals:
    Signal \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._Finished\: boolean := false;
    Signal \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0.return\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._Started\: boolean := false;
    Signal \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0.segmentSizeSize.parameter.In\: unsigned(7 downto 0) := to_unsigned(0, 8);
    -- System.UInt16 Lombiq.Unum.UnumHelper::SegmentSizeSizeToSegmentSize(System.Byte).0 declarations end


    -- System.Void Lombiq.Unum.UnumEnvironment::.ctor(System.Byte,System.Byte).0 declarations start
    -- State machine states:
    type \UnumEnvironment::.ctor(Byte,Byte).0._States\ is (
        \UnumEnvironment::.ctor(Byte,Byte).0._State_0\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_1\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_2\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_3\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_4\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_5\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_6\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_7\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_8\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_9\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_10\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_11\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_12\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_13\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_14\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_15\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_16\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_17\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_18\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_19\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_20\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_21\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_22\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_23\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_24\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_25\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_26\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_27\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_28\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_29\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_30\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_31\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_32\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_33\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_34\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_35\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_36\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_37\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_38\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_39\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_40\, 
        \UnumEnvironment::.ctor(Byte,Byte).0._State_41\);
    -- Signals:
    Signal \UnumEnvironment::.ctor(Byte,Byte).0._Finished\: boolean := false;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.this.parameter.Out\: \Lombiq.Unum.UnumEnvironment\;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.UnumHelper::SegmentSizeSizeToSegmentSize(Byte).segmentSizeSize.parameter.Out.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.UnumHelper::SegmentSizeSizeToSegmentSize(Byte)._Started.0\: boolean := false;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\: boolean := false;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\: boolean := false;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).this.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).index.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Started.0\: boolean := false;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).right.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\: boolean := false;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_BitwiseOr(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_BitwiseOr(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_BitwiseOr(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask).right.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\: boolean := false;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,UInt32).left.parameter.Out.0\: \Lombiq.Unum.BitMask\;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\: boolean := false;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0._Started\: boolean := false;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.this.parameter.In\: \Lombiq.Unum.UnumEnvironment\;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.exponentSizeSize.parameter.In\: unsigned(7 downto 0) := to_unsigned(0, 8);
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.fractionSizeSize.parameter.In\: unsigned(7 downto 0) := to_unsigned(0, 8);
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.UnumHelper::SegmentSizeSizeToSegmentSize(Byte)._Finished.0\: boolean := false;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.UnumHelper::SegmentSizeSizeToSegmentSize(Byte).return.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\: \Lombiq.Unum.BitMask\;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\: boolean := false;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Finished.0\: boolean := false;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).return.0\: \Lombiq.Unum.BitMask\;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\: boolean := false;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).return.0\: \Lombiq.Unum.BitMask\;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask).return.0\: \Lombiq.Unum.BitMask\;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_BitwiseOr(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_BitwiseOr(BitMask,BitMask).return.0\: \Lombiq.Unum.BitMask\;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\: boolean := false;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask).return.0\: \Lombiq.Unum.BitMask\;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\: boolean := false;
    Signal \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,UInt32).return.0\: \Lombiq.Unum.BitMask\;
    -- System.Void Lombiq.Unum.UnumEnvironment::.ctor(System.Byte,System.Byte).0 declarations end


    -- System.Void Hast::ExternalInvocationProxy() declarations start
    -- Signals:
    Signal \FinishedInternal\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory)._Finished.0\: boolean := false;
    -- System.Void Hast::ExternalInvocationProxy() declarations end


    -- \System.Void Hast::InternalInvocationProxy()._CommonDeclarations\ declarations start
    type \InternalInvocationProxy_boolean_Array\ is array (integer range <>) of boolean;
    type \Hast::InternalInvocationProxy()._RunningStates\ is (
        WaitingForStarted, 
        WaitingForFinished, 
        AfterFinished);
    -- \System.Void Hast::InternalInvocationProxy()._CommonDeclarations\ declarations end

begin 

    -- System.Void Hast.Samples.SampleAssembly.UnumCalculator::CalculateSumOfPowersofTwo(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine start
    \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._StateMachine\: process (\Clock\) 
        Variable \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\: \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._States\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_0\;
        Variable \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.environment\: \Lombiq.Unum.UnumEnvironment\;
        Variable \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.unum\: \Lombiq.Unum.Unum\;
        Variable \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.left\: \Lombiq.Unum.Unum\;
        Variable \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.num2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.array\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
        Variable \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.i\: signed(31 downto 0) := to_signed(0, 32);
        Variable \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.dataIn.0\: std_logic_vector(31 downto 0);
        Variable \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.return.0\: \Lombiq.Unum.UnumEnvironment\;
        Variable \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.0\: boolean := false;
        Variable \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.1\: boolean := false;
        Variable \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.return.1\: \Lombiq.Unum.Unum\;
        Variable \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.return.2\: \Lombiq.Unum.Unum\;
        Variable \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.return.3\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
        Variable \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.3\: boolean := false;
        Variable \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.4\: boolean := false;
        Variable \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.5\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._Finished\ <= false;
                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.UnumCalculator::EnvironmentFactory()._Started.0\ <= false;
                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32).value.parameter.Out.0\ <= to_signed(0, 32);
                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32)._Started.0\ <= false;
                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum)._Started.0\ <= false;
                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::FractionToUintArray()._Started.0\ <= false;
                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_0\;
                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.num\ := to_unsigned(0, 32);
                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.num2\ := to_signed(0, 32);
                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.array\ := (others => to_unsigned(0, 32));
                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.i\ := to_signed(0, 32);
                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.0\ := false;
                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.1\ := false;
                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.2\ := to_signed(0, 32);
                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.return.3\ := (others => to_unsigned(0, 32));
                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.3\ := false;
                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.4\ := false;
                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.5\ := to_signed(0, 32);
            else 
                case \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ is 
                    when \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._Started\ = true) then 
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._Started\ = true) then 
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._Finished\ <= true;
                        else 
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._Finished\ <= false;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_2\ => 
                        -- Begin SimpleMemory read.
                        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(to_signed(0, 32), 32);
                        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.SimpleMemory.ReadEnable\ <= true;
                        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_3\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\ReadsDone\ = true) then 
                            -- SimpleMemory read finished.
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.dataIn.0\ := \DataIn\;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.num\ := ConvertStdLogicVectorToUInt32(\UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.dataIn.0\);
                            -- Starting state machine invocation for the following method: Lombiq.Unum.UnumEnvironment Hast.Samples.SampleAssembly.UnumCalculator::EnvironmentFactory()
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.UnumCalculator::EnvironmentFactory()._Started.0\ <= true;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.UnumEnvironment Hast.Samples.SampleAssembly.UnumCalculator::EnvironmentFactory()
                        if (\UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.UnumCalculator::EnvironmentFactory()._Started.0\ = \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.UnumCalculator::EnvironmentFactory()._Finished.0\) then 
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.UnumCalculator::EnvironmentFactory()._Started.0\ <= false;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.return.0\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.UnumCalculator::EnvironmentFactory().return.0\;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.environment\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.return.0\;
                            -- Initializing record fields to their defaults.
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.unum\.\IsNull\ := false;
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.Int32)
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32).this.parameter.Out.0\ <= \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.unum\;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32).environment.parameter.Out.0\ <= \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.environment\;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32).value.parameter.Out.0\ <= to_signed(1, 32);
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32)._Started.0\ <= true;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.Int32)
                        if (\UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32)._Started.0\ = \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32)._Finished.0\) then 
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32)._Started.0\ <= false;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.unum\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32).this.parameter.In.0\;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.environment\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32).environment.parameter.In.0\;
                            -- Initializing record fields to their defaults.
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.left\.\IsNull\ := false;
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.Int32)
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32).this.parameter.Out.0\ <= \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.left\;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32).environment.parameter.Out.0\ <= \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.environment\;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32).value.parameter.Out.0\ <= to_signed(0, 32);
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32)._Started.0\ <= true;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_6\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.Int32)
                        if (\UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32)._Started.0\ = \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32)._Finished.0\) then 
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32)._Started.0\ <= false;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.left\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32).this.parameter.In.0\;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.environment\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32).environment.parameter.In.0\;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.num2\ := to_signed(1, 32);
                            -- Starting a while loop.
                            -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.0\ := resize(\UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.num2\, 64) <= signed((resize(\UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.num\, 64)));
                            if (\UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.0\) then 
                                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_7\;
                            else 
                                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_8\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_7\ => 
                        -- Repeated state of the while loop which was started in state \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_6\.
                        -- The while loop's condition:
                        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.1\ := resize(\UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.num2\, 64) <= signed((resize(\UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.num\, 64)));
                        if (\UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.1\) then 
                            -- Starting state machine invocation for the following method: Lombiq.Unum.Unum Lombiq.Unum.Unum::op_Addition(Lombiq.Unum.Unum,Lombiq.Unum.Unum)
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum).left.parameter.Out.0\ <= \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.left\;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum).right.parameter.Out.0\ <= \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.unum\;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum)._Started.0\ <= true;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_9\;
                        else 
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_8\ => 
                        -- State after the while loop which was started in state \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_6\.
                        -- Starting state machine invocation for the following method: System.UInt32[] Lombiq.Unum.Unum::FractionToUintArray()
                        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::FractionToUintArray().this.parameter.Out.0\ <= \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.left\;
                        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::FractionToUintArray()._Started.0\ <= true;
                        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_13\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_9\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.Unum Lombiq.Unum.Unum::op_Addition(Lombiq.Unum.Unum,Lombiq.Unum.Unum)
                        if (\UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum)._Started.0\ = \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum)._Finished.0\) then 
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum)._Started.0\ <= false;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.return.1\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum).return.0\;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.left\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.return.1\;
                            -- The last invocation for the target state machine just finished, so need to start the next one in a later state.
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_10\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_10\ => 
                        -- This state was just added to leave time for the invocation proxy to register that the previous invocation finished.
                        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_11\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_11\ => 
                        -- Starting state machine invocation for the following method: Lombiq.Unum.Unum Lombiq.Unum.Unum::op_Addition(Lombiq.Unum.Unum,Lombiq.Unum.Unum)
                        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum).left.parameter.Out.0\ <= \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.unum\;
                        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum).right.parameter.Out.0\ <= \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.unum\;
                        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum)._Started.0\ <= true;
                        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_12\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_12\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.Unum Lombiq.Unum.Unum::op_Addition(Lombiq.Unum.Unum,Lombiq.Unum.Unum)
                        if (\UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum)._Started.0\ = \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum)._Finished.0\) then 
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum)._Started.0\ <= false;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.return.2\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum).return.0\;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.unum\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.return.2\;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.2\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.num2\ + to_signed(1, 32);
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.num2\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.2\;
                            -- Returning to the repeated state of the while loop which was started in state \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_6\ if the loop wasn't exited with a state change.
                            if (\UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ = \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_12\) then 
                                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_7\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_13\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32[] Lombiq.Unum.Unum::FractionToUintArray()
                        if (\UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::FractionToUintArray()._Started.0\ = \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::FractionToUintArray()._Finished.0\) then 
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::FractionToUintArray()._Started.0\ <= false;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.return.3\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::FractionToUintArray().return.0\;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.array\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.return.3\;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.i\ := to_signed(0, 32);
                            -- Starting a while loop.
                            -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.3\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.i\ < to_signed(9, 32);
                            if (\UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.3\) then 
                                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_14\;
                            else 
                                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_15\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_14\ => 
                        -- Repeated state of the while loop which was started in state \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_13\.
                        -- The while loop's condition:
                        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.4\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.i\ < to_signed(9, 32);
                        if (\UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.4\) then 
                            -- Begin SimpleMemory write.
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.SimpleMemory.CellIndex\ <= resize(\UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.i\, 32);
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.SimpleMemory.WriteEnable\ <= true;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.SimpleMemory.DataOut\ <= ConvertUInt32ToStdLogicVector(\UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.array\(to_integer(\UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.i\)));
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_16\;
                        else 
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_15\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_15\ => 
                        -- State after the while loop which was started in state \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_13\.
                        \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_16\ => 
                        -- Waiting for the SimpleMemory operation to finish.
                        if (\WritesDone\ = true) then 
                            -- SimpleMemory write finished.
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.5\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.i\ + to_signed(1, 32);
                            \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.i\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.binaryOperationResult.5\;
                            -- Returning to the repeated state of the while loop which was started in state \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_13\ if the loop wasn't exited with a state change.
                            if (\UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ = \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_16\) then 
                                \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State\ := \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._State_14\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.Samples.SampleAssembly.UnumCalculator::CalculateSumOfPowersofTwo(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 state machine end


    -- Lombiq.Unum.UnumEnvironment Hast.Samples.SampleAssembly.UnumCalculator::EnvironmentFactory().0 state machine start
    \UnumCalculator::EnvironmentFactory().0._StateMachine\: process (\Clock\) 
        Variable \UnumCalculator::EnvironmentFactory().0._State\: \UnumCalculator::EnvironmentFactory().0._States\ := \UnumCalculator::EnvironmentFactory().0._State_0\;
        Variable \UnumCalculator::EnvironmentFactory().0.objectb022c2ea5fd837b49ebefe7712f46e723c82f78f2185697b6b6db16e6ca8c10d\: \Lombiq.Unum.UnumEnvironment\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \UnumCalculator::EnvironmentFactory().0._Finished\ <= false;
                \UnumCalculator::EnvironmentFactory().0.UnumEnvironment::.ctor(Byte,Byte).exponentSizeSize.parameter.Out.0\ <= to_unsigned(0, 8);
                \UnumCalculator::EnvironmentFactory().0.UnumEnvironment::.ctor(Byte,Byte).fractionSizeSize.parameter.Out.0\ <= to_unsigned(0, 8);
                \UnumCalculator::EnvironmentFactory().0.UnumEnvironment::.ctor(Byte,Byte)._Started.0\ <= false;
                \UnumCalculator::EnvironmentFactory().0._State\ := \UnumCalculator::EnvironmentFactory().0._State_0\;
            else 
                case \UnumCalculator::EnvironmentFactory().0._State\ is 
                    when \UnumCalculator::EnvironmentFactory().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\UnumCalculator::EnvironmentFactory().0._Started\ = true) then 
                            \UnumCalculator::EnvironmentFactory().0._State\ := \UnumCalculator::EnvironmentFactory().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumCalculator::EnvironmentFactory().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\UnumCalculator::EnvironmentFactory().0._Started\ = true) then 
                            \UnumCalculator::EnvironmentFactory().0._Finished\ <= true;
                        else 
                            \UnumCalculator::EnvironmentFactory().0._Finished\ <= false;
                            \UnumCalculator::EnvironmentFactory().0._State\ := \UnumCalculator::EnvironmentFactory().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumCalculator::EnvironmentFactory().0._State_2\ => 
                        -- Initializing record fields to their defaults.
                        \UnumCalculator::EnvironmentFactory().0.objectb022c2ea5fd837b49ebefe7712f46e723c82f78f2185697b6b6db16e6ca8c10d\.\IsNull\ := false;
                        \UnumCalculator::EnvironmentFactory().0.objectb022c2ea5fd837b49ebefe7712f46e723c82f78f2185697b6b6db16e6ca8c10d\.\ExponentSizeSize\ := to_unsigned(0, 8);
                        \UnumCalculator::EnvironmentFactory().0.objectb022c2ea5fd837b49ebefe7712f46e723c82f78f2185697b6b6db16e6ca8c10d\.\FractionSizeSize\ := to_unsigned(0, 8);
                        \UnumCalculator::EnvironmentFactory().0.objectb022c2ea5fd837b49ebefe7712f46e723c82f78f2185697b6b6db16e6ca8c10d\.\ExponentSizeMax\ := to_unsigned(0, 8);
                        \UnumCalculator::EnvironmentFactory().0.objectb022c2ea5fd837b49ebefe7712f46e723c82f78f2185697b6b6db16e6ca8c10d\.\FractionSizeMax\ := to_unsigned(0, 16);
                        \UnumCalculator::EnvironmentFactory().0.objectb022c2ea5fd837b49ebefe7712f46e723c82f78f2185697b6b6db16e6ca8c10d\.\UnumTagSize\ := to_unsigned(0, 8);
                        \UnumCalculator::EnvironmentFactory().0.objectb022c2ea5fd837b49ebefe7712f46e723c82f78f2185697b6b6db16e6ca8c10d\.\Size\ := to_unsigned(0, 16);
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.UnumEnvironment::.ctor(System.Byte,System.Byte)
                        \UnumCalculator::EnvironmentFactory().0.UnumEnvironment::.ctor(Byte,Byte).this.parameter.Out.0\ <= \UnumCalculator::EnvironmentFactory().0.objectb022c2ea5fd837b49ebefe7712f46e723c82f78f2185697b6b6db16e6ca8c10d\;
                        \UnumCalculator::EnvironmentFactory().0.UnumEnvironment::.ctor(Byte,Byte).exponentSizeSize.parameter.Out.0\ <= to_unsigned(4, 8);
                        \UnumCalculator::EnvironmentFactory().0.UnumEnvironment::.ctor(Byte,Byte).fractionSizeSize.parameter.Out.0\ <= to_unsigned(8, 8);
                        \UnumCalculator::EnvironmentFactory().0.UnumEnvironment::.ctor(Byte,Byte)._Started.0\ <= true;
                        \UnumCalculator::EnvironmentFactory().0._State\ := \UnumCalculator::EnvironmentFactory().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumCalculator::EnvironmentFactory().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.UnumEnvironment::.ctor(System.Byte,System.Byte)
                        if (\UnumCalculator::EnvironmentFactory().0.UnumEnvironment::.ctor(Byte,Byte)._Started.0\ = \UnumCalculator::EnvironmentFactory().0.UnumEnvironment::.ctor(Byte,Byte)._Finished.0\) then 
                            \UnumCalculator::EnvironmentFactory().0.UnumEnvironment::.ctor(Byte,Byte)._Started.0\ <= false;
                            \UnumCalculator::EnvironmentFactory().0.objectb022c2ea5fd837b49ebefe7712f46e723c82f78f2185697b6b6db16e6ca8c10d\ := \UnumCalculator::EnvironmentFactory().0.UnumEnvironment::.ctor(Byte,Byte).this.parameter.In.0\;
                            \UnumCalculator::EnvironmentFactory().0.return\ <= \UnumCalculator::EnvironmentFactory().0.objectb022c2ea5fd837b49ebefe7712f46e723c82f78f2185697b6b6db16e6ca8c10d\;
                            \UnumCalculator::EnvironmentFactory().0._State\ := \UnumCalculator::EnvironmentFactory().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.UnumEnvironment Hast.Samples.SampleAssembly.UnumCalculator::EnvironmentFactory().0 state machine end


    -- System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16).0 state machine start
    \BitMask::.ctor(UInt32[],UInt16).0._StateMachine\: process (\Clock\) 
        Variable \BitMask::.ctor(UInt32[],UInt16).0._State\: \BitMask::.ctor(UInt32[],UInt16).0._States\ := \BitMask::.ctor(UInt32[],UInt16).0._State_0\;
        Variable \BitMask::.ctor(UInt32[],UInt16).0.this\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::.ctor(UInt32[],UInt16).0.segments\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
        Variable \BitMask::.ctor(UInt32[],UInt16).0.size\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::.ctor(UInt32[],UInt16).0.num\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::.ctor(UInt32[],UInt16).0.flag\: boolean := false;
        Variable \BitMask::.ctor(UInt32[],UInt16).0.array\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
        Variable \BitMask::.ctor(UInt32[],UInt16).0.conditionalc3a7314574e5cf5b60b9437fa75a8e8b23417040c5c46d12edec97fe2eb66018\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.0\: boolean := false;
        Variable \BitMask::.ctor(UInt32[],UInt16).0.conditional93d0384e1e256fd728e80c772ac32f7836cc8471edbcd4a0afb4c8bc9bb86ec2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.1\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::.ctor(UInt32[],UInt16).0.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.2\: boolean := false;
        Variable \BitMask::.ctor(UInt32[],UInt16).0.conditionalb63e6b911b0b9623cc84e1b95d8ef143c98867889a1ec5a3ac70836cafbf43ac\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.3\: boolean := false;
        Variable \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.4\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.5\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.6\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \BitMask::.ctor(UInt32[],UInt16).0._Finished\ <= false;
                \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.Out\ <= (others => to_unsigned(0, 32));
                \BitMask::.ctor(UInt32[],UInt16).0._State\ := \BitMask::.ctor(UInt32[],UInt16).0._State_0\;
                \BitMask::.ctor(UInt32[],UInt16).0.segments\ := (others => to_unsigned(0, 32));
                \BitMask::.ctor(UInt32[],UInt16).0.size\ := to_unsigned(0, 16);
                \BitMask::.ctor(UInt32[],UInt16).0.num\ := to_unsigned(0, 16);
                \BitMask::.ctor(UInt32[],UInt16).0.flag\ := false;
                \BitMask::.ctor(UInt32[],UInt16).0.array\ := (others => to_unsigned(0, 32));
                \BitMask::.ctor(UInt32[],UInt16).0.conditionalc3a7314574e5cf5b60b9437fa75a8e8b23417040c5c46d12edec97fe2eb66018\ := to_unsigned(0, 16);
                \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.0\ := false;
                \BitMask::.ctor(UInt32[],UInt16).0.conditional93d0384e1e256fd728e80c772ac32f7836cc8471edbcd4a0afb4c8bc9bb86ec2\ := to_signed(0, 32);
                \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.1\ := to_unsigned(0, 16);
                \BitMask::.ctor(UInt32[],UInt16).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.2\ := false;
                \BitMask::.ctor(UInt32[],UInt16).0.conditionalb63e6b911b0b9623cc84e1b95d8ef143c98867889a1ec5a3ac70836cafbf43ac\ := to_unsigned(0, 16);
                \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.3\ := false;
                \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.4\ := to_signed(0, 32);
                \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.5\ := to_unsigned(0, 16);
                \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.6\ := false;
            else 
                case \BitMask::.ctor(UInt32[],UInt16).0._State\ is 
                    when \BitMask::.ctor(UInt32[],UInt16).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\BitMask::.ctor(UInt32[],UInt16).0._Started\ = true) then 
                            \BitMask::.ctor(UInt32[],UInt16).0._State\ := \BitMask::.ctor(UInt32[],UInt16).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::.ctor(UInt32[],UInt16).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\BitMask::.ctor(UInt32[],UInt16).0._Started\ = true) then 
                            \BitMask::.ctor(UInt32[],UInt16).0._Finished\ <= true;
                        else 
                            \BitMask::.ctor(UInt32[],UInt16).0._Finished\ <= false;
                            \BitMask::.ctor(UInt32[],UInt16).0._State\ := \BitMask::.ctor(UInt32[],UInt16).0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.Out\ <= \BitMask::.ctor(UInt32[],UInt16).0.this\;
                        \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.Out\ <= \BitMask::.ctor(UInt32[],UInt16).0.segments\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::.ctor(UInt32[],UInt16).0._State_2\ => 
                        \BitMask::.ctor(UInt32[],UInt16).0.this\ := \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.In\;
                        \BitMask::.ctor(UInt32[],UInt16).0.segments\ := \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.In\;
                        \BitMask::.ctor(UInt32[],UInt16).0.size\ := \BitMask::.ctor(UInt32[],UInt16).0.size.parameter.In\;
                        \BitMask::.ctor(UInt32[],UInt16).0.num\ := to_unsigned(288, 16);
                        \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.0\ := \BitMask::.ctor(UInt32[],UInt16).0.size\ < to_unsigned(288, 16);

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::.ctor(UInt32[],UInt16).0._State_4\ and ends in state \BitMask::.ctor(UInt32[],UInt16).0._State_4\.
                        --     * The false branch starts in state \BitMask::.ctor(UInt32[],UInt16).0._State_5\ and ends in state \BitMask::.ctor(UInt32[],UInt16).0._State_5\.
                        --     * Execution after either branch will continue in the following state: \BitMask::.ctor(UInt32[],UInt16).0._State_3\.

                        if (\BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.0\) then 
                            \BitMask::.ctor(UInt32[],UInt16).0._State\ := \BitMask::.ctor(UInt32[],UInt16).0._State_4\;
                        else 
                            \BitMask::.ctor(UInt32[],UInt16).0._State\ := \BitMask::.ctor(UInt32[],UInt16).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::.ctor(UInt32[],UInt16).0._State_3\ => 
                        -- State after the if-else which was started in state \BitMask::.ctor(UInt32[],UInt16).0._State_2\.
                        \BitMask::.ctor(UInt32[],UInt16).0.this\.\Size\ := \BitMask::.ctor(UInt32[],UInt16).0.conditionalc3a7314574e5cf5b60b9437fa75a8e8b23417040c5c46d12edec97fe2eb66018\;
                        \BitMask::.ctor(UInt32[],UInt16).0._State\ := \BitMask::.ctor(UInt32[],UInt16).0._State_6\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::.ctor(UInt32[],UInt16).0._State_4\ => 
                        -- True branch of the if-else started in state \BitMask::.ctor(UInt32[],UInt16).0._State_2\.
                        \BitMask::.ctor(UInt32[],UInt16).0.conditionalc3a7314574e5cf5b60b9437fa75a8e8b23417040c5c46d12edec97fe2eb66018\ := to_unsigned(288, 16);
                        -- Going to the state after the if-else which was started in state \BitMask::.ctor(UInt32[],UInt16).0._State_2\.
                        if (\BitMask::.ctor(UInt32[],UInt16).0._State\ = \BitMask::.ctor(UInt32[],UInt16).0._State_4\) then 
                            \BitMask::.ctor(UInt32[],UInt16).0._State\ := \BitMask::.ctor(UInt32[],UInt16).0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::.ctor(UInt32[],UInt16).0._State_5\ => 
                        -- False branch of the if-else started in state \BitMask::.ctor(UInt32[],UInt16).0._State_2\.
                        \BitMask::.ctor(UInt32[],UInt16).0.conditionalc3a7314574e5cf5b60b9437fa75a8e8b23417040c5c46d12edec97fe2eb66018\ := \BitMask::.ctor(UInt32[],UInt16).0.size\;
                        -- Going to the state after the if-else which was started in state \BitMask::.ctor(UInt32[],UInt16).0._State_2\.
                        if (\BitMask::.ctor(UInt32[],UInt16).0._State\ = \BitMask::.ctor(UInt32[],UInt16).0._State_5\) then 
                            \BitMask::.ctor(UInt32[],UInt16).0._State\ := \BitMask::.ctor(UInt32[],UInt16).0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::.ctor(UInt32[],UInt16).0._State_6\ => 
                        -- Waiting for the result to appear in \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.1\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\BitMask::.ctor(UInt32[],UInt16).0.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \BitMask::.ctor(UInt32[],UInt16).0._State\ := \BitMask::.ctor(UInt32[],UInt16).0._State_7\;
                            \BitMask::.ctor(UInt32[],UInt16).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \BitMask::.ctor(UInt32[],UInt16).0.clockCyclesWaitedForBinaryOperationResult.0\ := \BitMask::.ctor(UInt32[],UInt16).0.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.1\ := \BitMask::.ctor(UInt32[],UInt16).0.size\ mod to_unsigned(32, 16);
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \BitMask::.ctor(UInt32[],UInt16).0._State_7\ => 
                        \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.2\ := \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.1\ = to_unsigned(0, 16);

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::.ctor(UInt32[],UInt16).0._State_9\ and ends in state \BitMask::.ctor(UInt32[],UInt16).0._State_9\.
                        --     * The false branch starts in state \BitMask::.ctor(UInt32[],UInt16).0._State_10\ and ends in state \BitMask::.ctor(UInt32[],UInt16).0._State_10\.
                        --     * Execution after either branch will continue in the following state: \BitMask::.ctor(UInt32[],UInt16).0._State_8\.

                        if (\BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.2\) then 
                            \BitMask::.ctor(UInt32[],UInt16).0._State\ := \BitMask::.ctor(UInt32[],UInt16).0._State_9\;
                        else 
                            \BitMask::.ctor(UInt32[],UInt16).0._State\ := \BitMask::.ctor(UInt32[],UInt16).0._State_10\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::.ctor(UInt32[],UInt16).0._State_8\ => 
                        -- State after the if-else which was started in state \BitMask::.ctor(UInt32[],UInt16).0._State_7\.
                        \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.3\ := \BitMask::.ctor(UInt32[],UInt16).0.size\ > to_unsigned(288, 16);

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::.ctor(UInt32[],UInt16).0._State_12\ and ends in state \BitMask::.ctor(UInt32[],UInt16).0._State_12\.
                        --     * The false branch starts in state \BitMask::.ctor(UInt32[],UInt16).0._State_13\ and ends in state \BitMask::.ctor(UInt32[],UInt16).0._State_13\.
                        --     * Execution after either branch will continue in the following state: \BitMask::.ctor(UInt32[],UInt16).0._State_11\.

                        if (\BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.3\) then 
                            \BitMask::.ctor(UInt32[],UInt16).0._State\ := \BitMask::.ctor(UInt32[],UInt16).0._State_12\;
                        else 
                            \BitMask::.ctor(UInt32[],UInt16).0._State\ := \BitMask::.ctor(UInt32[],UInt16).0._State_13\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::.ctor(UInt32[],UInt16).0._State_9\ => 
                        -- True branch of the if-else started in state \BitMask::.ctor(UInt32[],UInt16).0._State_7\.
                        \BitMask::.ctor(UInt32[],UInt16).0.conditional93d0384e1e256fd728e80c772ac32f7836cc8471edbcd4a0afb4c8bc9bb86ec2\ := to_signed(0, 32);
                        -- Going to the state after the if-else which was started in state \BitMask::.ctor(UInt32[],UInt16).0._State_7\.
                        if (\BitMask::.ctor(UInt32[],UInt16).0._State\ = \BitMask::.ctor(UInt32[],UInt16).0._State_9\) then 
                            \BitMask::.ctor(UInt32[],UInt16).0._State\ := \BitMask::.ctor(UInt32[],UInt16).0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::.ctor(UInt32[],UInt16).0._State_10\ => 
                        -- False branch of the if-else started in state \BitMask::.ctor(UInt32[],UInt16).0._State_7\.
                        \BitMask::.ctor(UInt32[],UInt16).0.conditional93d0384e1e256fd728e80c772ac32f7836cc8471edbcd4a0afb4c8bc9bb86ec2\ := to_signed(1, 32);
                        -- Going to the state after the if-else which was started in state \BitMask::.ctor(UInt32[],UInt16).0._State_7\.
                        if (\BitMask::.ctor(UInt32[],UInt16).0._State\ = \BitMask::.ctor(UInt32[],UInt16).0._State_10\) then 
                            \BitMask::.ctor(UInt32[],UInt16).0._State\ := \BitMask::.ctor(UInt32[],UInt16).0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::.ctor(UInt32[],UInt16).0._State_11\ => 
                        -- State after the if-else which was started in state \BitMask::.ctor(UInt32[],UInt16).0._State_8\.
                        \BitMask::.ctor(UInt32[],UInt16).0.this\.\SegmentCount\ := \BitMask::.ctor(UInt32[],UInt16).0.conditionalb63e6b911b0b9623cc84e1b95d8ef143c98867889a1ec5a3ac70836cafbf43ac\;
                        \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.6\ := resize(signed(\BitMask::.ctor(UInt32[],UInt16).0.this\.\SegmentCount\), 32) > to_signed(9, 32);
                        \BitMask::.ctor(UInt32[],UInt16).0.flag\ := \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.6\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::.ctor(UInt32[],UInt16).0._State_15\ and ends in state \BitMask::.ctor(UInt32[],UInt16).0._State_15\.
                        --     * The false branch starts in state \BitMask::.ctor(UInt32[],UInt16).0._State_16\ and ends in state \BitMask::.ctor(UInt32[],UInt16).0._State_16\.
                        --     * Execution after either branch will continue in the following state: \BitMask::.ctor(UInt32[],UInt16).0._State_14\.

                        if (\BitMask::.ctor(UInt32[],UInt16).0.flag\) then 
                            \BitMask::.ctor(UInt32[],UInt16).0._State\ := \BitMask::.ctor(UInt32[],UInt16).0._State_15\;
                        else 
                            \BitMask::.ctor(UInt32[],UInt16).0._State\ := \BitMask::.ctor(UInt32[],UInt16).0._State_16\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::.ctor(UInt32[],UInt16).0._State_12\ => 
                        -- True branch of the if-else started in state \BitMask::.ctor(UInt32[],UInt16).0._State_8\.
                        \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.4\ := resize(signed(shift_right(\BitMask::.ctor(UInt32[],UInt16).0.size\, to_integer(to_signed(5, 32)))), 32);
                        \BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.5\ := resize(unsigned(\BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.4\ + \BitMask::.ctor(UInt32[],UInt16).0.conditional93d0384e1e256fd728e80c772ac32f7836cc8471edbcd4a0afb4c8bc9bb86ec2\), 16);
                        \BitMask::.ctor(UInt32[],UInt16).0.conditionalb63e6b911b0b9623cc84e1b95d8ef143c98867889a1ec5a3ac70836cafbf43ac\ := (\BitMask::.ctor(UInt32[],UInt16).0.binaryOperationResult.5\);
                        -- Going to the state after the if-else which was started in state \BitMask::.ctor(UInt32[],UInt16).0._State_8\.
                        if (\BitMask::.ctor(UInt32[],UInt16).0._State\ = \BitMask::.ctor(UInt32[],UInt16).0._State_12\) then 
                            \BitMask::.ctor(UInt32[],UInt16).0._State\ := \BitMask::.ctor(UInt32[],UInt16).0._State_11\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \BitMask::.ctor(UInt32[],UInt16).0._State_13\ => 
                        -- False branch of the if-else started in state \BitMask::.ctor(UInt32[],UInt16).0._State_8\.
                        \BitMask::.ctor(UInt32[],UInt16).0.conditionalb63e6b911b0b9623cc84e1b95d8ef143c98867889a1ec5a3ac70836cafbf43ac\ := to_unsigned(9, 16);
                        -- Going to the state after the if-else which was started in state \BitMask::.ctor(UInt32[],UInt16).0._State_8\.
                        if (\BitMask::.ctor(UInt32[],UInt16).0._State\ = \BitMask::.ctor(UInt32[],UInt16).0._State_13\) then 
                            \BitMask::.ctor(UInt32[],UInt16).0._State\ := \BitMask::.ctor(UInt32[],UInt16).0._State_11\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::.ctor(UInt32[],UInt16).0._State_14\ => 
                        -- State after the if-else which was started in state \BitMask::.ctor(UInt32[],UInt16).0._State_11\.
                        \BitMask::.ctor(UInt32[],UInt16).0._State\ := \BitMask::.ctor(UInt32[],UInt16).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::.ctor(UInt32[],UInt16).0._State_15\ => 
                        -- True branch of the if-else started in state \BitMask::.ctor(UInt32[],UInt16).0._State_11\.
                        \BitMask::.ctor(UInt32[],UInt16).0.array\ := (others => to_unsigned(0, 32));
                        \BitMask::.ctor(UInt32[],UInt16).0.array\ := \BitMask::.ctor(UInt32[],UInt16).0.segments\(0 to 8);
                        \BitMask::.ctor(UInt32[],UInt16).0.this\.\Segments\ := \BitMask::.ctor(UInt32[],UInt16).0.array\;
                        -- Going to the state after the if-else which was started in state \BitMask::.ctor(UInt32[],UInt16).0._State_11\.
                        if (\BitMask::.ctor(UInt32[],UInt16).0._State\ = \BitMask::.ctor(UInt32[],UInt16).0._State_15\) then 
                            \BitMask::.ctor(UInt32[],UInt16).0._State\ := \BitMask::.ctor(UInt32[],UInt16).0._State_14\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::.ctor(UInt32[],UInt16).0._State_16\ => 
                        -- False branch of the if-else started in state \BitMask::.ctor(UInt32[],UInt16).0._State_11\.
                        \BitMask::.ctor(UInt32[],UInt16).0.this\.\Segments\ := \BitMask::.ctor(UInt32[],UInt16).0.segments\;
                        -- Going to the state after the if-else which was started in state \BitMask::.ctor(UInt32[],UInt16).0._State_11\.
                        if (\BitMask::.ctor(UInt32[],UInt16).0._State\ = \BitMask::.ctor(UInt32[],UInt16).0._State_16\) then 
                            \BitMask::.ctor(UInt32[],UInt16).0._State\ := \BitMask::.ctor(UInt32[],UInt16).0._State_14\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16).0 state machine end


    -- System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean).0 state machine start
    \BitMask::.ctor(UInt16,Boolean).0._StateMachine\: process (\Clock\) 
        Variable \BitMask::.ctor(UInt16,Boolean).0._State\: \BitMask::.ctor(UInt16,Boolean).0._States\ := \BitMask::.ctor(UInt16,Boolean).0._State_0\;
        Variable \BitMask::.ctor(UInt16,Boolean).0.this\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::.ctor(UInt16,Boolean).0.size\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::.ctor(UInt16,Boolean).0.allOne\: boolean := false;
        Variable \BitMask::.ctor(UInt16,Boolean).0.num\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::.ctor(UInt16,Boolean).0.array\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
        Variable \BitMask::.ctor(UInt16,Boolean).0.num2\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::.ctor(UInt16,Boolean).0.binaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::.ctor(UInt16,Boolean).0.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::.ctor(UInt16,Boolean).0.conditional48feffe0202fc0c0df2cb980716aa7461c00997856cf3b8aeb212a7a22e7f468\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::.ctor(UInt16,Boolean).0.binaryOperationResult.1\: boolean := false;
        Variable \BitMask::.ctor(UInt16,Boolean).0.binaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::.ctor(UInt16,Boolean).0.binaryOperationResult.3\: unsigned(15 downto 0) := to_unsigned(0, 16);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \BitMask::.ctor(UInt16,Boolean).0._Finished\ <= false;
                \BitMask::.ctor(UInt16,Boolean).0._State\ := \BitMask::.ctor(UInt16,Boolean).0._State_0\;
                \BitMask::.ctor(UInt16,Boolean).0.size\ := to_unsigned(0, 16);
                \BitMask::.ctor(UInt16,Boolean).0.allOne\ := false;
                \BitMask::.ctor(UInt16,Boolean).0.num\ := to_signed(0, 32);
                \BitMask::.ctor(UInt16,Boolean).0.array\ := (others => to_unsigned(0, 32));
                \BitMask::.ctor(UInt16,Boolean).0.num2\ := to_unsigned(0, 16);
                \BitMask::.ctor(UInt16,Boolean).0.binaryOperationResult.0\ := to_signed(0, 32);
                \BitMask::.ctor(UInt16,Boolean).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                \BitMask::.ctor(UInt16,Boolean).0.conditional48feffe0202fc0c0df2cb980716aa7461c00997856cf3b8aeb212a7a22e7f468\ := to_signed(0, 32);
                \BitMask::.ctor(UInt16,Boolean).0.binaryOperationResult.1\ := false;
                \BitMask::.ctor(UInt16,Boolean).0.binaryOperationResult.2\ := to_signed(0, 32);
                \BitMask::.ctor(UInt16,Boolean).0.binaryOperationResult.3\ := to_unsigned(0, 16);
            else 
                case \BitMask::.ctor(UInt16,Boolean).0._State\ is 
                    when \BitMask::.ctor(UInt16,Boolean).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\BitMask::.ctor(UInt16,Boolean).0._Started\ = true) then 
                            \BitMask::.ctor(UInt16,Boolean).0._State\ := \BitMask::.ctor(UInt16,Boolean).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::.ctor(UInt16,Boolean).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\BitMask::.ctor(UInt16,Boolean).0._Started\ = true) then 
                            \BitMask::.ctor(UInt16,Boolean).0._Finished\ <= true;
                        else 
                            \BitMask::.ctor(UInt16,Boolean).0._Finished\ <= false;
                            \BitMask::.ctor(UInt16,Boolean).0._State\ := \BitMask::.ctor(UInt16,Boolean).0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \BitMask::.ctor(UInt16,Boolean).0.this.parameter.Out\ <= \BitMask::.ctor(UInt16,Boolean).0.this\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::.ctor(UInt16,Boolean).0._State_2\ => 
                        \BitMask::.ctor(UInt16,Boolean).0.this\ := \BitMask::.ctor(UInt16,Boolean).0.this.parameter.In\;
                        \BitMask::.ctor(UInt16,Boolean).0.size\ := \BitMask::.ctor(UInt16,Boolean).0.size.parameter.In\;
                        \BitMask::.ctor(UInt16,Boolean).0.allOne\ := \BitMask::.ctor(UInt16,Boolean).0.allOne.parameter.In\;
                        \BitMask::.ctor(UInt16,Boolean).0._State\ := \BitMask::.ctor(UInt16,Boolean).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::.ctor(UInt16,Boolean).0._State_3\ => 
                        -- Waiting for the result to appear in \BitMask::.ctor(UInt16,Boolean).0.binaryOperationResult.0\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\BitMask::.ctor(UInt16,Boolean).0.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \BitMask::.ctor(UInt16,Boolean).0._State\ := \BitMask::.ctor(UInt16,Boolean).0._State_4\;
                            \BitMask::.ctor(UInt16,Boolean).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \BitMask::.ctor(UInt16,Boolean).0.clockCyclesWaitedForBinaryOperationResult.0\ := \BitMask::.ctor(UInt16,Boolean).0.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        \BitMask::.ctor(UInt16,Boolean).0.binaryOperationResult.0\ := resize(signed(\BitMask::.ctor(UInt16,Boolean).0.size\ mod to_unsigned(32, 16)), 32);
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \BitMask::.ctor(UInt16,Boolean).0._State_4\ => 
                        \BitMask::.ctor(UInt16,Boolean).0.num\ := (\BitMask::.ctor(UInt16,Boolean).0.binaryOperationResult.0\);
                        \BitMask::.ctor(UInt16,Boolean).0.binaryOperationResult.1\ := \BitMask::.ctor(UInt16,Boolean).0.num\ = to_signed(0, 32);

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::.ctor(UInt16,Boolean).0._State_6\ and ends in state \BitMask::.ctor(UInt16,Boolean).0._State_6\.
                        --     * The false branch starts in state \BitMask::.ctor(UInt16,Boolean).0._State_7\ and ends in state \BitMask::.ctor(UInt16,Boolean).0._State_7\.
                        --     * Execution after either branch will continue in the following state: \BitMask::.ctor(UInt16,Boolean).0._State_5\.

                        if (\BitMask::.ctor(UInt16,Boolean).0.binaryOperationResult.1\) then 
                            \BitMask::.ctor(UInt16,Boolean).0._State\ := \BitMask::.ctor(UInt16,Boolean).0._State_6\;
                        else 
                            \BitMask::.ctor(UInt16,Boolean).0._State\ := \BitMask::.ctor(UInt16,Boolean).0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::.ctor(UInt16,Boolean).0._State_5\ => 
                        -- State after the if-else which was started in state \BitMask::.ctor(UInt16,Boolean).0._State_4\.
                        \BitMask::.ctor(UInt16,Boolean).0.binaryOperationResult.2\ := resize(signed(shift_right(\BitMask::.ctor(UInt16,Boolean).0.size\, to_integer(to_signed(5, 32)))), 32);
                        \BitMask::.ctor(UInt16,Boolean).0.binaryOperationResult.3\ := resize(unsigned(\BitMask::.ctor(UInt16,Boolean).0.binaryOperationResult.2\ + \BitMask::.ctor(UInt16,Boolean).0.conditional48feffe0202fc0c0df2cb980716aa7461c00997856cf3b8aeb212a7a22e7f468\), 16);
                        \BitMask::.ctor(UInt16,Boolean).0.this\.\SegmentCount\ := (\BitMask::.ctor(UInt16,Boolean).0.binaryOperationResult.3\);
                        \BitMask::.ctor(UInt16,Boolean).0.this\.\Size\ := \BitMask::.ctor(UInt16,Boolean).0.size\;
                        \BitMask::.ctor(UInt16,Boolean).0.array\ := (others => to_unsigned(0, 32));
                        \BitMask::.ctor(UInt16,Boolean).0.this\.\Segments\ := \BitMask::.ctor(UInt16,Boolean).0.array\;
                        \BitMask::.ctor(UInt16,Boolean).0._State\ := \BitMask::.ctor(UInt16,Boolean).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \BitMask::.ctor(UInt16,Boolean).0._State_6\ => 
                        -- True branch of the if-else started in state \BitMask::.ctor(UInt16,Boolean).0._State_4\.
                        \BitMask::.ctor(UInt16,Boolean).0.conditional48feffe0202fc0c0df2cb980716aa7461c00997856cf3b8aeb212a7a22e7f468\ := to_signed(0, 32);
                        -- Going to the state after the if-else which was started in state \BitMask::.ctor(UInt16,Boolean).0._State_4\.
                        if (\BitMask::.ctor(UInt16,Boolean).0._State\ = \BitMask::.ctor(UInt16,Boolean).0._State_6\) then 
                            \BitMask::.ctor(UInt16,Boolean).0._State\ := \BitMask::.ctor(UInt16,Boolean).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::.ctor(UInt16,Boolean).0._State_7\ => 
                        -- False branch of the if-else started in state \BitMask::.ctor(UInt16,Boolean).0._State_4\.
                        \BitMask::.ctor(UInt16,Boolean).0.conditional48feffe0202fc0c0df2cb980716aa7461c00997856cf3b8aeb212a7a22e7f468\ := to_signed(1, 32);
                        -- Going to the state after the if-else which was started in state \BitMask::.ctor(UInt16,Boolean).0._State_4\.
                        if (\BitMask::.ctor(UInt16,Boolean).0._State\ = \BitMask::.ctor(UInt16,Boolean).0._State_7\) then 
                            \BitMask::.ctor(UInt16,Boolean).0._State\ := \BitMask::.ctor(UInt16,Boolean).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean).0 state machine end


    -- System.Void Lombiq.Unum.BitMask::.ctor(Lombiq.Unum.BitMask).0 state machine start
    \BitMask::.ctor(BitMask).0._StateMachine\: process (\Clock\) 
        Variable \BitMask::.ctor(BitMask).0._State\: \BitMask::.ctor(BitMask).0._States\ := \BitMask::.ctor(BitMask).0._State_0\;
        Variable \BitMask::.ctor(BitMask).0.this\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::.ctor(BitMask).0.source\: \Lombiq.Unum.BitMask\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \BitMask::.ctor(BitMask).0._Finished\ <= false;
                \BitMask::.ctor(BitMask).0._State\ := \BitMask::.ctor(BitMask).0._State_0\;
            else 
                case \BitMask::.ctor(BitMask).0._State\ is 
                    when \BitMask::.ctor(BitMask).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\BitMask::.ctor(BitMask).0._Started\ = true) then 
                            \BitMask::.ctor(BitMask).0._State\ := \BitMask::.ctor(BitMask).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::.ctor(BitMask).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\BitMask::.ctor(BitMask).0._Started\ = true) then 
                            \BitMask::.ctor(BitMask).0._Finished\ <= true;
                        else 
                            \BitMask::.ctor(BitMask).0._Finished\ <= false;
                            \BitMask::.ctor(BitMask).0._State\ := \BitMask::.ctor(BitMask).0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \BitMask::.ctor(BitMask).0.this.parameter.Out\ <= \BitMask::.ctor(BitMask).0.this\;
                        \BitMask::.ctor(BitMask).0.source.parameter.Out\ <= \BitMask::.ctor(BitMask).0.source\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::.ctor(BitMask).0._State_2\ => 
                        \BitMask::.ctor(BitMask).0.this\ := \BitMask::.ctor(BitMask).0.this.parameter.In\;
                        \BitMask::.ctor(BitMask).0.source\ := \BitMask::.ctor(BitMask).0.source.parameter.In\;
                        \BitMask::.ctor(BitMask).0.this\.\Size\ := \BitMask::.ctor(BitMask).0.source\.\Size\;
                        \BitMask::.ctor(BitMask).0.this\.\SegmentCount\ := \BitMask::.ctor(BitMask).0.source\.\SegmentCount\;
                        \BitMask::.ctor(BitMask).0.this\.\Segments\ := \BitMask::.ctor(BitMask).0.source\.\Segments\;
                        \BitMask::.ctor(BitMask).0._State\ := \BitMask::.ctor(BitMask).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Lombiq.Unum.BitMask::.ctor(Lombiq.Unum.BitMask).0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::FromImmutableArray(System.UInt32[],System.UInt16).0 state machine start
    \BitMask::FromImmutableArray(UInt32[],UInt16).0._StateMachine\: process (\Clock\) 
        Variable \BitMask::FromImmutableArray(UInt32[],UInt16).0._State\: \BitMask::FromImmutableArray(UInt32[],UInt16).0._States\ := \BitMask::FromImmutableArray(UInt32[],UInt16).0._State_0\;
        Variable \BitMask::FromImmutableArray(UInt32[],UInt16).0.segments\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
        Variable \BitMask::FromImmutableArray(UInt32[],UInt16).0.size\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::FromImmutableArray(UInt32[],UInt16).0.array\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
        Variable \BitMask::FromImmutableArray(UInt32[],UInt16).0.object2fe313ea47a5c88e5364ea75f59651d95bb221efab0dda850bcb112321cfbdac\: \Lombiq.Unum.BitMask\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \BitMask::FromImmutableArray(UInt32[],UInt16).0._Finished\ <= false;
                \BitMask::FromImmutableArray(UInt32[],UInt16).0.segments.parameter.Out\ <= (others => to_unsigned(0, 32));
                \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 32));
                \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                \BitMask::FromImmutableArray(UInt32[],UInt16).0._State\ := \BitMask::FromImmutableArray(UInt32[],UInt16).0._State_0\;
                \BitMask::FromImmutableArray(UInt32[],UInt16).0.segments\ := (others => to_unsigned(0, 32));
                \BitMask::FromImmutableArray(UInt32[],UInt16).0.size\ := to_unsigned(0, 16);
                \BitMask::FromImmutableArray(UInt32[],UInt16).0.array\ := (others => to_unsigned(0, 32));
            else 
                case \BitMask::FromImmutableArray(UInt32[],UInt16).0._State\ is 
                    when \BitMask::FromImmutableArray(UInt32[],UInt16).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\BitMask::FromImmutableArray(UInt32[],UInt16).0._Started\ = true) then 
                            \BitMask::FromImmutableArray(UInt32[],UInt16).0._State\ := \BitMask::FromImmutableArray(UInt32[],UInt16).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::FromImmutableArray(UInt32[],UInt16).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\BitMask::FromImmutableArray(UInt32[],UInt16).0._Started\ = true) then 
                            \BitMask::FromImmutableArray(UInt32[],UInt16).0._Finished\ <= true;
                        else 
                            \BitMask::FromImmutableArray(UInt32[],UInt16).0._Finished\ <= false;
                            \BitMask::FromImmutableArray(UInt32[],UInt16).0._State\ := \BitMask::FromImmutableArray(UInt32[],UInt16).0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \BitMask::FromImmutableArray(UInt32[],UInt16).0.segments.parameter.Out\ <= \BitMask::FromImmutableArray(UInt32[],UInt16).0.segments\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::FromImmutableArray(UInt32[],UInt16).0._State_2\ => 
                        \BitMask::FromImmutableArray(UInt32[],UInt16).0.segments\ := \BitMask::FromImmutableArray(UInt32[],UInt16).0.segments.parameter.In\;
                        \BitMask::FromImmutableArray(UInt32[],UInt16).0.size\ := \BitMask::FromImmutableArray(UInt32[],UInt16).0.size.parameter.In\;
                        \BitMask::FromImmutableArray(UInt32[],UInt16).0.array\ := (others => to_unsigned(0, 32));
                        \BitMask::FromImmutableArray(UInt32[],UInt16).0.array\ := \BitMask::FromImmutableArray(UInt32[],UInt16).0.segments\(0 to 8);
                        -- Initializing record fields to their defaults.
                        \BitMask::FromImmutableArray(UInt32[],UInt16).0.object2fe313ea47a5c88e5364ea75f59651d95bb221efab0dda850bcb112321cfbdac\.\IsNull\ := false;
                        \BitMask::FromImmutableArray(UInt32[],UInt16).0.object2fe313ea47a5c88e5364ea75f59651d95bb221efab0dda850bcb112321cfbdac\.\Size\ := to_unsigned(0, 16);
                        \BitMask::FromImmutableArray(UInt32[],UInt16).0.object2fe313ea47a5c88e5364ea75f59651d95bb221efab0dda850bcb112321cfbdac\.\SegmentCount\ := to_unsigned(0, 16);
                        \BitMask::FromImmutableArray(UInt32[],UInt16).0.object2fe313ea47a5c88e5364ea75f59651d95bb221efab0dda850bcb112321cfbdac\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\ <= \BitMask::FromImmutableArray(UInt32[],UInt16).0.object2fe313ea47a5c88e5364ea75f59651d95bb221efab0dda850bcb112321cfbdac\;
                        \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\ <= \BitMask::FromImmutableArray(UInt32[],UInt16).0.array\;
                        \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= \BitMask::FromImmutableArray(UInt32[],UInt16).0.size\;
                        \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= true;
                        \BitMask::FromImmutableArray(UInt32[],UInt16).0._State\ := \BitMask::FromImmutableArray(UInt32[],UInt16).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::FromImmutableArray(UInt32[],UInt16).0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        if (\BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\) then 
                            \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                            \BitMask::FromImmutableArray(UInt32[],UInt16).0.object2fe313ea47a5c88e5364ea75f59651d95bb221efab0dda850bcb112321cfbdac\ := \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\;
                            \BitMask::FromImmutableArray(UInt32[],UInt16).0.array\ := \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\;
                            \BitMask::FromImmutableArray(UInt32[],UInt16).0.return\ <= \BitMask::FromImmutableArray(UInt32[],UInt16).0.object2fe313ea47a5c88e5364ea75f59651d95bb221efab0dda850bcb112321cfbdac\;
                            \BitMask::FromImmutableArray(UInt32[],UInt16).0._State\ := \BitMask::FromImmutableArray(UInt32[],UInt16).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::FromImmutableArray(System.UInt32[],System.UInt16).0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetOne(System.UInt16).0 state machine start
    \BitMask::SetOne(UInt16).0._StateMachine\: process (\Clock\) 
        Variable \BitMask::SetOne(UInt16).0._State\: \BitMask::SetOne(UInt16).0._States\ := \BitMask::SetOne(UInt16).0._State_0\;
        Variable \BitMask::SetOne(UInt16).0.this\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::SetOne(UInt16).0.index\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::SetOne(UInt16).0.flag\: boolean := false;
        Variable \BitMask::SetOne(UInt16).0.result\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::SetOne(UInt16).0.num\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::SetOne(UInt16).0.index2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::SetOne(UInt16).0.flag2\: boolean := false;
        Variable \BitMask::SetOne(UInt16).0.binaryOperationResult.0\: boolean := false;
        Variable \BitMask::SetOne(UInt16).0.binaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::SetOne(UInt16).0.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::SetOne(UInt16).0.binaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::SetOne(UInt16).0.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::SetOne(UInt16).0.binaryOperationResult.4\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::SetOne(UInt16).0.clockCyclesWaitedForBinaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::SetOne(UInt16).0.binaryOperationResult.5\: boolean := false;
        Variable \BitMask::SetOne(UInt16).0.arraya674cb90f8197922d5e1ac95ff9cb374a98401cf0158bcfad208496fd1c9c68c\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
        Variable \BitMask::SetOne(UInt16).0.binaryOperationResult.6\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::SetOne(UInt16).0.binaryOperationResult.7\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::SetOne(UInt16).0.return.0\: \Lombiq.Unum.BitMask\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \BitMask::SetOne(UInt16).0._Finished\ <= false;
                \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask)._Started.0\ <= false;
                \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 32));
                \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Started.0\ <= false;
                \BitMask::SetOne(UInt16).0._State\ := \BitMask::SetOne(UInt16).0._State_0\;
                \BitMask::SetOne(UInt16).0.index\ := to_unsigned(0, 16);
                \BitMask::SetOne(UInt16).0.flag\ := false;
                \BitMask::SetOne(UInt16).0.num\ := to_signed(0, 32);
                \BitMask::SetOne(UInt16).0.index2\ := to_signed(0, 32);
                \BitMask::SetOne(UInt16).0.flag2\ := false;
                \BitMask::SetOne(UInt16).0.binaryOperationResult.0\ := false;
                \BitMask::SetOne(UInt16).0.binaryOperationResult.1\ := to_signed(0, 32);
                \BitMask::SetOne(UInt16).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                \BitMask::SetOne(UInt16).0.binaryOperationResult.2\ := to_signed(0, 32);
                \BitMask::SetOne(UInt16).0.binaryOperationResult.3\ := to_unsigned(0, 32);
                \BitMask::SetOne(UInt16).0.binaryOperationResult.4\ := to_unsigned(0, 32);
                \BitMask::SetOne(UInt16).0.clockCyclesWaitedForBinaryOperationResult.1\ := to_signed(0, 32);
                \BitMask::SetOne(UInt16).0.binaryOperationResult.5\ := false;
                \BitMask::SetOne(UInt16).0.arraya674cb90f8197922d5e1ac95ff9cb374a98401cf0158bcfad208496fd1c9c68c\ := (others => to_unsigned(0, 32));
                \BitMask::SetOne(UInt16).0.binaryOperationResult.6\ := to_unsigned(0, 32);
                \BitMask::SetOne(UInt16).0.binaryOperationResult.7\ := to_unsigned(0, 32);
            else 
                case \BitMask::SetOne(UInt16).0._State\ is 
                    when \BitMask::SetOne(UInt16).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\BitMask::SetOne(UInt16).0._Started\ = true) then 
                            \BitMask::SetOne(UInt16).0._State\ := \BitMask::SetOne(UInt16).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::SetOne(UInt16).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\BitMask::SetOne(UInt16).0._Started\ = true) then 
                            \BitMask::SetOne(UInt16).0._Finished\ <= true;
                        else 
                            \BitMask::SetOne(UInt16).0._Finished\ <= false;
                            \BitMask::SetOne(UInt16).0._State\ := \BitMask::SetOne(UInt16).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::SetOne(UInt16).0._State_2\ => 
                        \BitMask::SetOne(UInt16).0.this\ := \BitMask::SetOne(UInt16).0.this.parameter.In\;
                        \BitMask::SetOne(UInt16).0.index\ := \BitMask::SetOne(UInt16).0.index.parameter.In\;
                        \BitMask::SetOne(UInt16).0.binaryOperationResult.0\ := \BitMask::SetOne(UInt16).0.index\ > \BitMask::SetOne(UInt16).0.this\.\Size\;
                        \BitMask::SetOne(UInt16).0.flag\ := \BitMask::SetOne(UInt16).0.binaryOperationResult.0\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::SetOne(UInt16).0._State_4\ and ends in state \BitMask::SetOne(UInt16).0._State_5\.
                        --     * The false branch starts in state \BitMask::SetOne(UInt16).0._State_6\ and ends in state \BitMask::SetOne(UInt16).0._State_11\.
                        --     * Execution after either branch will continue in the following state: \BitMask::SetOne(UInt16).0._State_3\.

                        if (\BitMask::SetOne(UInt16).0.flag\) then 
                            \BitMask::SetOne(UInt16).0._State\ := \BitMask::SetOne(UInt16).0._State_4\;
                        else 
                            \BitMask::SetOne(UInt16).0._State\ := \BitMask::SetOne(UInt16).0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::SetOne(UInt16).0._State_3\ => 
                        -- State after the if-else which was started in state \BitMask::SetOne(UInt16).0._State_2\.
                        \BitMask::SetOne(UInt16).0.return\ <= \BitMask::SetOne(UInt16).0.result\;
                        \BitMask::SetOne(UInt16).0._State\ := \BitMask::SetOne(UInt16).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::SetOne(UInt16).0._State_4\ => 
                        -- True branch of the if-else started in state \BitMask::SetOne(UInt16).0._State_2\.
                        -- Initializing record fields to their defaults.
                        \BitMask::SetOne(UInt16).0.result\.\IsNull\ := false;
                        \BitMask::SetOne(UInt16).0.result\.\Size\ := to_unsigned(0, 16);
                        \BitMask::SetOne(UInt16).0.result\.\SegmentCount\ := to_unsigned(0, 16);
                        \BitMask::SetOne(UInt16).0.result\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(Lombiq.Unum.BitMask)
                        \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask).this.parameter.Out.0\ <= \BitMask::SetOne(UInt16).0.result\;
                        \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask).source.parameter.Out.0\ <= \BitMask::SetOne(UInt16).0.this\;
                        \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask)._Started.0\ <= true;
                        \BitMask::SetOne(UInt16).0._State\ := \BitMask::SetOne(UInt16).0._State_5\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::SetOne(UInt16).0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(Lombiq.Unum.BitMask)
                        if (\BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask)._Started.0\ = \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask)._Finished.0\) then 
                            \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask)._Started.0\ <= false;
                            \BitMask::SetOne(UInt16).0.result\ := \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask).this.parameter.In.0\;
                            \BitMask::SetOne(UInt16).0.this\ := \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask).source.parameter.In.0\;
                            -- Going to the state after the if-else which was started in state \BitMask::SetOne(UInt16).0._State_2\.
                            if (\BitMask::SetOne(UInt16).0._State\ = \BitMask::SetOne(UInt16).0._State_5\) then 
                                \BitMask::SetOne(UInt16).0._State\ := \BitMask::SetOne(UInt16).0._State_3\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::SetOne(UInt16).0._State_6\ => 
                        -- False branch of the if-else started in state \BitMask::SetOne(UInt16).0._State_2\.
                        \BitMask::SetOne(UInt16).0._State\ := \BitMask::SetOne(UInt16).0._State_7\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::SetOne(UInt16).0._State_7\ => 
                        -- Waiting for the result to appear in \BitMask::SetOne(UInt16).0.binaryOperationResult.1\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\BitMask::SetOne(UInt16).0.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \BitMask::SetOne(UInt16).0._State\ := \BitMask::SetOne(UInt16).0._State_8\;
                            \BitMask::SetOne(UInt16).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \BitMask::SetOne(UInt16).0.clockCyclesWaitedForBinaryOperationResult.0\ := \BitMask::SetOne(UInt16).0.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        \BitMask::SetOne(UInt16).0.binaryOperationResult.1\ := resize(signed(\BitMask::SetOne(UInt16).0.index\ mod to_unsigned(32, 16)), 32);
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \BitMask::SetOne(UInt16).0._State_8\ => 
                        \BitMask::SetOne(UInt16).0.num\ := (\BitMask::SetOne(UInt16).0.binaryOperationResult.1\);
                        \BitMask::SetOne(UInt16).0.binaryOperationResult.2\ := resize(signed(shift_right(\BitMask::SetOne(UInt16).0.index\, to_integer(to_signed(5, 32)))), 32);
                        \BitMask::SetOne(UInt16).0.index2\ := \BitMask::SetOne(UInt16).0.binaryOperationResult.2\;
                        \BitMask::SetOne(UInt16).0.binaryOperationResult.3\ := shift_right(\BitMask::SetOne(UInt16).0.this\.\Segments\(to_integer(\BitMask::SetOne(UInt16).0.index2\)), to_integer(unsigned(\BitMask::SetOne(UInt16).0.num\)));
                        \BitMask::SetOne(UInt16).0._State\ := \BitMask::SetOne(UInt16).0._State_9\;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \BitMask::SetOne(UInt16).0._State_9\ => 
                        -- Waiting for the result to appear in \BitMask::SetOne(UInt16).0.binaryOperationResult.4\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\BitMask::SetOne(UInt16).0.clockCyclesWaitedForBinaryOperationResult.1\ >= to_signed(7, 32)) then 
                            \BitMask::SetOne(UInt16).0._State\ := \BitMask::SetOne(UInt16).0._State_10\;
                            \BitMask::SetOne(UInt16).0.clockCyclesWaitedForBinaryOperationResult.1\ := to_signed(0, 32);
                        else 
                            \BitMask::SetOne(UInt16).0.clockCyclesWaitedForBinaryOperationResult.1\ := \BitMask::SetOne(UInt16).0.clockCyclesWaitedForBinaryOperationResult.1\ + to_signed(1, 32);
                        end if;
                        \BitMask::SetOne(UInt16).0.binaryOperationResult.4\ := \BitMask::SetOne(UInt16).0.binaryOperationResult.3\ mod to_unsigned(2, 32);
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \BitMask::SetOne(UInt16).0._State_10\ => 
                        \BitMask::SetOne(UInt16).0.binaryOperationResult.5\ := \BitMask::SetOne(UInt16).0.binaryOperationResult.4\ = to_unsigned(0, 32);
                        \BitMask::SetOne(UInt16).0.flag2\ := \BitMask::SetOne(UInt16).0.binaryOperationResult.5\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::SetOne(UInt16).0._State_12\ and ends in state \BitMask::SetOne(UInt16).0._State_13\.
                        --     * The false branch starts in state \BitMask::SetOne(UInt16).0._State_14\ and ends in state \BitMask::SetOne(UInt16).0._State_15\.
                        --     * Execution after either branch will continue in the following state: \BitMask::SetOne(UInt16).0._State_11\.

                        if (\BitMask::SetOne(UInt16).0.flag2\) then 
                            \BitMask::SetOne(UInt16).0._State\ := \BitMask::SetOne(UInt16).0._State_12\;
                        else 
                            \BitMask::SetOne(UInt16).0._State\ := \BitMask::SetOne(UInt16).0._State_14\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::SetOne(UInt16).0._State_11\ => 
                        -- State after the if-else which was started in state \BitMask::SetOne(UInt16).0._State_10\.
                        -- Going to the state after the if-else which was started in state \BitMask::SetOne(UInt16).0._State_2\.
                        if (\BitMask::SetOne(UInt16).0._State\ = \BitMask::SetOne(UInt16).0._State_11\) then 
                            \BitMask::SetOne(UInt16).0._State\ := \BitMask::SetOne(UInt16).0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::SetOne(UInt16).0._State_12\ => 
                        -- True branch of the if-else started in state \BitMask::SetOne(UInt16).0._State_10\.
                        \BitMask::SetOne(UInt16).0.arraya674cb90f8197922d5e1ac95ff9cb374a98401cf0158bcfad208496fd1c9c68c\ := (others => to_unsigned(0, 32));
                        \BitMask::SetOne(UInt16).0.arraya674cb90f8197922d5e1ac95ff9cb374a98401cf0158bcfad208496fd1c9c68c\ := \BitMask::SetOne(UInt16).0.this\.\Segments\(0 to 8);
                        \BitMask::SetOne(UInt16).0.binaryOperationResult.6\ := shift_left(to_unsigned(1, 32), to_integer(\BitMask::SetOne(UInt16).0.num\));
                        \BitMask::SetOne(UInt16).0.binaryOperationResult.7\ := \BitMask::SetOne(UInt16).0.this\.\Segments\(to_integer(\BitMask::SetOne(UInt16).0.index2\)) or \BitMask::SetOne(UInt16).0.binaryOperationResult.6\;
                        \BitMask::SetOne(UInt16).0.arraya674cb90f8197922d5e1ac95ff9cb374a98401cf0158bcfad208496fd1c9c68c\(to_integer(\BitMask::SetOne(UInt16).0.index2\)) := \BitMask::SetOne(UInt16).0.binaryOperationResult.7\;
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::FromImmutableArray(System.UInt32[],System.UInt16)
                        \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).segments.parameter.Out.0\ <= \BitMask::SetOne(UInt16).0.arraya674cb90f8197922d5e1ac95ff9cb374a98401cf0158bcfad208496fd1c9c68c\;
                        \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).size.parameter.Out.0\ <= \BitMask::SetOne(UInt16).0.this\.\Size\;
                        \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Started.0\ <= true;
                        \BitMask::SetOne(UInt16).0._State\ := \BitMask::SetOne(UInt16).0._State_13\;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \BitMask::SetOne(UInt16).0._State_13\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::FromImmutableArray(System.UInt32[],System.UInt16)
                        if (\BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Started.0\ = \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Finished.0\) then 
                            \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Started.0\ <= false;
                            \BitMask::SetOne(UInt16).0.return.0\ := \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).return.0\;
                            \BitMask::SetOne(UInt16).0.arraya674cb90f8197922d5e1ac95ff9cb374a98401cf0158bcfad208496fd1c9c68c\ := \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).segments.parameter.In.0\;
                            \BitMask::SetOne(UInt16).0.result\ := \BitMask::SetOne(UInt16).0.return.0\;
                            -- Going to the state after the if-else which was started in state \BitMask::SetOne(UInt16).0._State_10\.
                            if (\BitMask::SetOne(UInt16).0._State\ = \BitMask::SetOne(UInt16).0._State_13\) then 
                                \BitMask::SetOne(UInt16).0._State\ := \BitMask::SetOne(UInt16).0._State_11\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::SetOne(UInt16).0._State_14\ => 
                        -- False branch of the if-else started in state \BitMask::SetOne(UInt16).0._State_10\.
                        -- Initializing record fields to their defaults.
                        \BitMask::SetOne(UInt16).0.result\.\IsNull\ := false;
                        \BitMask::SetOne(UInt16).0.result\.\Size\ := to_unsigned(0, 16);
                        \BitMask::SetOne(UInt16).0.result\.\SegmentCount\ := to_unsigned(0, 16);
                        \BitMask::SetOne(UInt16).0.result\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(Lombiq.Unum.BitMask)
                        \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask).this.parameter.Out.0\ <= \BitMask::SetOne(UInt16).0.result\;
                        \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask).source.parameter.Out.0\ <= \BitMask::SetOne(UInt16).0.this\;
                        \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask)._Started.0\ <= true;
                        \BitMask::SetOne(UInt16).0._State\ := \BitMask::SetOne(UInt16).0._State_15\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::SetOne(UInt16).0._State_15\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(Lombiq.Unum.BitMask)
                        if (\BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask)._Started.0\ = \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask)._Finished.0\) then 
                            \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask)._Started.0\ <= false;
                            \BitMask::SetOne(UInt16).0.result\ := \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask).this.parameter.In.0\;
                            \BitMask::SetOne(UInt16).0.this\ := \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask).source.parameter.In.0\;
                            -- Going to the state after the if-else which was started in state \BitMask::SetOne(UInt16).0._State_10\.
                            if (\BitMask::SetOne(UInt16).0._State\ = \BitMask::SetOne(UInt16).0._State_15\) then 
                                \BitMask::SetOne(UInt16).0._State\ := \BitMask::SetOne(UInt16).0._State_11\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetOne(System.UInt16).0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetZero(System.UInt16).0 state machine start
    \BitMask::SetZero(UInt16).0._StateMachine\: process (\Clock\) 
        Variable \BitMask::SetZero(UInt16).0._State\: \BitMask::SetZero(UInt16).0._States\ := \BitMask::SetZero(UInt16).0._State_0\;
        Variable \BitMask::SetZero(UInt16).0.this\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::SetZero(UInt16).0.index\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::SetZero(UInt16).0.flag\: boolean := false;
        Variable \BitMask::SetZero(UInt16).0.result\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::SetZero(UInt16).0.num\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::SetZero(UInt16).0.index2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::SetZero(UInt16).0.flag2\: boolean := false;
        Variable \BitMask::SetZero(UInt16).0.binaryOperationResult.0\: boolean := false;
        Variable \BitMask::SetZero(UInt16).0.binaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::SetZero(UInt16).0.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::SetZero(UInt16).0.binaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::SetZero(UInt16).0.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::SetZero(UInt16).0.binaryOperationResult.4\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::SetZero(UInt16).0.clockCyclesWaitedForBinaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::SetZero(UInt16).0.binaryOperationResult.5\: boolean := false;
        Variable \BitMask::SetZero(UInt16).0.array3d06f98f2942194f65130a81f3bd43f7302c3ca1bd92e1393a1cf0bfd23292c5\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
        Variable \BitMask::SetZero(UInt16).0.binaryOperationResult.6\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::SetZero(UInt16).0.binaryOperationResult.7\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::SetZero(UInt16).0.return.0\: \Lombiq.Unum.BitMask\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \BitMask::SetZero(UInt16).0._Finished\ <= false;
                \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask)._Started.0\ <= false;
                \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 32));
                \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Started.0\ <= false;
                \BitMask::SetZero(UInt16).0._State\ := \BitMask::SetZero(UInt16).0._State_0\;
                \BitMask::SetZero(UInt16).0.index\ := to_unsigned(0, 16);
                \BitMask::SetZero(UInt16).0.flag\ := false;
                \BitMask::SetZero(UInt16).0.num\ := to_signed(0, 32);
                \BitMask::SetZero(UInt16).0.index2\ := to_signed(0, 32);
                \BitMask::SetZero(UInt16).0.flag2\ := false;
                \BitMask::SetZero(UInt16).0.binaryOperationResult.0\ := false;
                \BitMask::SetZero(UInt16).0.binaryOperationResult.1\ := to_signed(0, 32);
                \BitMask::SetZero(UInt16).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                \BitMask::SetZero(UInt16).0.binaryOperationResult.2\ := to_signed(0, 32);
                \BitMask::SetZero(UInt16).0.binaryOperationResult.3\ := to_unsigned(0, 32);
                \BitMask::SetZero(UInt16).0.binaryOperationResult.4\ := to_unsigned(0, 32);
                \BitMask::SetZero(UInt16).0.clockCyclesWaitedForBinaryOperationResult.1\ := to_signed(0, 32);
                \BitMask::SetZero(UInt16).0.binaryOperationResult.5\ := false;
                \BitMask::SetZero(UInt16).0.array3d06f98f2942194f65130a81f3bd43f7302c3ca1bd92e1393a1cf0bfd23292c5\ := (others => to_unsigned(0, 32));
                \BitMask::SetZero(UInt16).0.binaryOperationResult.6\ := to_unsigned(0, 32);
                \BitMask::SetZero(UInt16).0.binaryOperationResult.7\ := to_unsigned(0, 32);
            else 
                case \BitMask::SetZero(UInt16).0._State\ is 
                    when \BitMask::SetZero(UInt16).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\BitMask::SetZero(UInt16).0._Started\ = true) then 
                            \BitMask::SetZero(UInt16).0._State\ := \BitMask::SetZero(UInt16).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::SetZero(UInt16).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\BitMask::SetZero(UInt16).0._Started\ = true) then 
                            \BitMask::SetZero(UInt16).0._Finished\ <= true;
                        else 
                            \BitMask::SetZero(UInt16).0._Finished\ <= false;
                            \BitMask::SetZero(UInt16).0._State\ := \BitMask::SetZero(UInt16).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::SetZero(UInt16).0._State_2\ => 
                        \BitMask::SetZero(UInt16).0.this\ := \BitMask::SetZero(UInt16).0.this.parameter.In\;
                        \BitMask::SetZero(UInt16).0.index\ := \BitMask::SetZero(UInt16).0.index.parameter.In\;
                        \BitMask::SetZero(UInt16).0.binaryOperationResult.0\ := \BitMask::SetZero(UInt16).0.index\ > \BitMask::SetZero(UInt16).0.this\.\Size\;
                        \BitMask::SetZero(UInt16).0.flag\ := \BitMask::SetZero(UInt16).0.binaryOperationResult.0\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::SetZero(UInt16).0._State_4\ and ends in state \BitMask::SetZero(UInt16).0._State_5\.
                        --     * The false branch starts in state \BitMask::SetZero(UInt16).0._State_6\ and ends in state \BitMask::SetZero(UInt16).0._State_11\.
                        --     * Execution after either branch will continue in the following state: \BitMask::SetZero(UInt16).0._State_3\.

                        if (\BitMask::SetZero(UInt16).0.flag\) then 
                            \BitMask::SetZero(UInt16).0._State\ := \BitMask::SetZero(UInt16).0._State_4\;
                        else 
                            \BitMask::SetZero(UInt16).0._State\ := \BitMask::SetZero(UInt16).0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::SetZero(UInt16).0._State_3\ => 
                        -- State after the if-else which was started in state \BitMask::SetZero(UInt16).0._State_2\.
                        \BitMask::SetZero(UInt16).0.return\ <= \BitMask::SetZero(UInt16).0.result\;
                        \BitMask::SetZero(UInt16).0._State\ := \BitMask::SetZero(UInt16).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::SetZero(UInt16).0._State_4\ => 
                        -- True branch of the if-else started in state \BitMask::SetZero(UInt16).0._State_2\.
                        -- Initializing record fields to their defaults.
                        \BitMask::SetZero(UInt16).0.result\.\IsNull\ := false;
                        \BitMask::SetZero(UInt16).0.result\.\Size\ := to_unsigned(0, 16);
                        \BitMask::SetZero(UInt16).0.result\.\SegmentCount\ := to_unsigned(0, 16);
                        \BitMask::SetZero(UInt16).0.result\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(Lombiq.Unum.BitMask)
                        \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask).this.parameter.Out.0\ <= \BitMask::SetZero(UInt16).0.result\;
                        \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask).source.parameter.Out.0\ <= \BitMask::SetZero(UInt16).0.this\;
                        \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask)._Started.0\ <= true;
                        \BitMask::SetZero(UInt16).0._State\ := \BitMask::SetZero(UInt16).0._State_5\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::SetZero(UInt16).0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(Lombiq.Unum.BitMask)
                        if (\BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask)._Started.0\ = \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask)._Finished.0\) then 
                            \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask)._Started.0\ <= false;
                            \BitMask::SetZero(UInt16).0.result\ := \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask).this.parameter.In.0\;
                            \BitMask::SetZero(UInt16).0.this\ := \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask).source.parameter.In.0\;
                            -- Going to the state after the if-else which was started in state \BitMask::SetZero(UInt16).0._State_2\.
                            if (\BitMask::SetZero(UInt16).0._State\ = \BitMask::SetZero(UInt16).0._State_5\) then 
                                \BitMask::SetZero(UInt16).0._State\ := \BitMask::SetZero(UInt16).0._State_3\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::SetZero(UInt16).0._State_6\ => 
                        -- False branch of the if-else started in state \BitMask::SetZero(UInt16).0._State_2\.
                        \BitMask::SetZero(UInt16).0._State\ := \BitMask::SetZero(UInt16).0._State_7\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::SetZero(UInt16).0._State_7\ => 
                        -- Waiting for the result to appear in \BitMask::SetZero(UInt16).0.binaryOperationResult.1\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\BitMask::SetZero(UInt16).0.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \BitMask::SetZero(UInt16).0._State\ := \BitMask::SetZero(UInt16).0._State_8\;
                            \BitMask::SetZero(UInt16).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \BitMask::SetZero(UInt16).0.clockCyclesWaitedForBinaryOperationResult.0\ := \BitMask::SetZero(UInt16).0.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        \BitMask::SetZero(UInt16).0.binaryOperationResult.1\ := resize(signed(\BitMask::SetZero(UInt16).0.index\ mod to_unsigned(32, 16)), 32);
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \BitMask::SetZero(UInt16).0._State_8\ => 
                        \BitMask::SetZero(UInt16).0.num\ := (\BitMask::SetZero(UInt16).0.binaryOperationResult.1\);
                        \BitMask::SetZero(UInt16).0.binaryOperationResult.2\ := resize(signed(shift_right(\BitMask::SetZero(UInt16).0.index\, to_integer(to_signed(5, 32)))), 32);
                        \BitMask::SetZero(UInt16).0.index2\ := \BitMask::SetZero(UInt16).0.binaryOperationResult.2\;
                        \BitMask::SetZero(UInt16).0.binaryOperationResult.3\ := shift_right(\BitMask::SetZero(UInt16).0.this\.\Segments\(to_integer(\BitMask::SetZero(UInt16).0.index2\)), to_integer(unsigned(\BitMask::SetZero(UInt16).0.num\)));
                        \BitMask::SetZero(UInt16).0._State\ := \BitMask::SetZero(UInt16).0._State_9\;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \BitMask::SetZero(UInt16).0._State_9\ => 
                        -- Waiting for the result to appear in \BitMask::SetZero(UInt16).0.binaryOperationResult.4\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\BitMask::SetZero(UInt16).0.clockCyclesWaitedForBinaryOperationResult.1\ >= to_signed(7, 32)) then 
                            \BitMask::SetZero(UInt16).0._State\ := \BitMask::SetZero(UInt16).0._State_10\;
                            \BitMask::SetZero(UInt16).0.clockCyclesWaitedForBinaryOperationResult.1\ := to_signed(0, 32);
                        else 
                            \BitMask::SetZero(UInt16).0.clockCyclesWaitedForBinaryOperationResult.1\ := \BitMask::SetZero(UInt16).0.clockCyclesWaitedForBinaryOperationResult.1\ + to_signed(1, 32);
                        end if;
                        \BitMask::SetZero(UInt16).0.binaryOperationResult.4\ := \BitMask::SetZero(UInt16).0.binaryOperationResult.3\ mod to_unsigned(2, 32);
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \BitMask::SetZero(UInt16).0._State_10\ => 
                        \BitMask::SetZero(UInt16).0.binaryOperationResult.5\ := \BitMask::SetZero(UInt16).0.binaryOperationResult.4\ = to_unsigned(1, 32);
                        \BitMask::SetZero(UInt16).0.flag2\ := \BitMask::SetZero(UInt16).0.binaryOperationResult.5\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::SetZero(UInt16).0._State_12\ and ends in state \BitMask::SetZero(UInt16).0._State_13\.
                        --     * The false branch starts in state \BitMask::SetZero(UInt16).0._State_14\ and ends in state \BitMask::SetZero(UInt16).0._State_15\.
                        --     * Execution after either branch will continue in the following state: \BitMask::SetZero(UInt16).0._State_11\.

                        if (\BitMask::SetZero(UInt16).0.flag2\) then 
                            \BitMask::SetZero(UInt16).0._State\ := \BitMask::SetZero(UInt16).0._State_12\;
                        else 
                            \BitMask::SetZero(UInt16).0._State\ := \BitMask::SetZero(UInt16).0._State_14\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::SetZero(UInt16).0._State_11\ => 
                        -- State after the if-else which was started in state \BitMask::SetZero(UInt16).0._State_10\.
                        -- Going to the state after the if-else which was started in state \BitMask::SetZero(UInt16).0._State_2\.
                        if (\BitMask::SetZero(UInt16).0._State\ = \BitMask::SetZero(UInt16).0._State_11\) then 
                            \BitMask::SetZero(UInt16).0._State\ := \BitMask::SetZero(UInt16).0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::SetZero(UInt16).0._State_12\ => 
                        -- True branch of the if-else started in state \BitMask::SetZero(UInt16).0._State_10\.
                        \BitMask::SetZero(UInt16).0.array3d06f98f2942194f65130a81f3bd43f7302c3ca1bd92e1393a1cf0bfd23292c5\ := (others => to_unsigned(0, 32));
                        \BitMask::SetZero(UInt16).0.array3d06f98f2942194f65130a81f3bd43f7302c3ca1bd92e1393a1cf0bfd23292c5\ := \BitMask::SetZero(UInt16).0.this\.\Segments\(0 to 8);
                        \BitMask::SetZero(UInt16).0.binaryOperationResult.6\ := shift_left(to_unsigned(1, 32), to_integer(\BitMask::SetZero(UInt16).0.num\));
                        \BitMask::SetZero(UInt16).0.binaryOperationResult.7\ := \BitMask::SetZero(UInt16).0.this\.\Segments\(to_integer(\BitMask::SetZero(UInt16).0.index2\)) and not(\BitMask::SetZero(UInt16).0.binaryOperationResult.6\);
                        \BitMask::SetZero(UInt16).0.array3d06f98f2942194f65130a81f3bd43f7302c3ca1bd92e1393a1cf0bfd23292c5\(to_integer(\BitMask::SetZero(UInt16).0.index2\)) := \BitMask::SetZero(UInt16).0.binaryOperationResult.7\;
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::FromImmutableArray(System.UInt32[],System.UInt16)
                        \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).segments.parameter.Out.0\ <= \BitMask::SetZero(UInt16).0.array3d06f98f2942194f65130a81f3bd43f7302c3ca1bd92e1393a1cf0bfd23292c5\;
                        \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).size.parameter.Out.0\ <= \BitMask::SetZero(UInt16).0.this\.\Size\;
                        \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Started.0\ <= true;
                        \BitMask::SetZero(UInt16).0._State\ := \BitMask::SetZero(UInt16).0._State_13\;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \BitMask::SetZero(UInt16).0._State_13\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::FromImmutableArray(System.UInt32[],System.UInt16)
                        if (\BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Started.0\ = \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Finished.0\) then 
                            \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Started.0\ <= false;
                            \BitMask::SetZero(UInt16).0.return.0\ := \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).return.0\;
                            \BitMask::SetZero(UInt16).0.array3d06f98f2942194f65130a81f3bd43f7302c3ca1bd92e1393a1cf0bfd23292c5\ := \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).segments.parameter.In.0\;
                            \BitMask::SetZero(UInt16).0.result\ := \BitMask::SetZero(UInt16).0.return.0\;
                            -- Going to the state after the if-else which was started in state \BitMask::SetZero(UInt16).0._State_10\.
                            if (\BitMask::SetZero(UInt16).0._State\ = \BitMask::SetZero(UInt16).0._State_13\) then 
                                \BitMask::SetZero(UInt16).0._State\ := \BitMask::SetZero(UInt16).0._State_11\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::SetZero(UInt16).0._State_14\ => 
                        -- False branch of the if-else started in state \BitMask::SetZero(UInt16).0._State_10\.
                        -- Initializing record fields to their defaults.
                        \BitMask::SetZero(UInt16).0.result\.\IsNull\ := false;
                        \BitMask::SetZero(UInt16).0.result\.\Size\ := to_unsigned(0, 16);
                        \BitMask::SetZero(UInt16).0.result\.\SegmentCount\ := to_unsigned(0, 16);
                        \BitMask::SetZero(UInt16).0.result\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(Lombiq.Unum.BitMask)
                        \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask).this.parameter.Out.0\ <= \BitMask::SetZero(UInt16).0.result\;
                        \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask).source.parameter.Out.0\ <= \BitMask::SetZero(UInt16).0.this\;
                        \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask)._Started.0\ <= true;
                        \BitMask::SetZero(UInt16).0._State\ := \BitMask::SetZero(UInt16).0._State_15\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::SetZero(UInt16).0._State_15\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(Lombiq.Unum.BitMask)
                        if (\BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask)._Started.0\ = \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask)._Finished.0\) then 
                            \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask)._Started.0\ <= false;
                            \BitMask::SetZero(UInt16).0.result\ := \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask).this.parameter.In.0\;
                            \BitMask::SetZero(UInt16).0.this\ := \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask).source.parameter.In.0\;
                            -- Going to the state after the if-else which was started in state \BitMask::SetZero(UInt16).0._State_10\.
                            if (\BitMask::SetZero(UInt16).0._State\ = \BitMask::SetZero(UInt16).0._State_15\) then 
                                \BitMask::SetZero(UInt16).0._State\ := \BitMask::SetZero(UInt16).0._State_11\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetZero(System.UInt16).0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::ShiftOutLeastSignificantZeros().0 state machine start
    \BitMask::ShiftOutLeastSignificantZeros().0._StateMachine\: process (\Clock\) 
        Variable \BitMask::ShiftOutLeastSignificantZeros().0._State\: \BitMask::ShiftOutLeastSignificantZeros().0._States\ := \BitMask::ShiftOutLeastSignificantZeros().0._State_0\;
        Variable \BitMask::ShiftOutLeastSignificantZeros().0.this\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::ShiftOutLeastSignificantZeros().0.leastSignificantOnePosition\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::ShiftOutLeastSignificantZeros().0.bitMask\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::ShiftOutLeastSignificantZeros().0.flag\: boolean := false;
        Variable \BitMask::ShiftOutLeastSignificantZeros().0.result\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::ShiftOutLeastSignificantZeros().0.return.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::ShiftOutLeastSignificantZeros().0.binaryOperationResult.0\: boolean := false;
        Variable \BitMask::ShiftOutLeastSignificantZeros().0.binaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::ShiftOutLeastSignificantZeros().0.return.1\: \Lombiq.Unum.BitMask\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \BitMask::ShiftOutLeastSignificantZeros().0._Finished\ <= false;
                \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::GetLeastSignificantOnePosition()._Started.0\ <= false;
                \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask)._Started.0\ <= false;
                \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::op_RightShift(BitMask,Int32).right.parameter.Out.0\ <= to_signed(0, 32);
                \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ <= false;
                \BitMask::ShiftOutLeastSignificantZeros().0._State\ := \BitMask::ShiftOutLeastSignificantZeros().0._State_0\;
                \BitMask::ShiftOutLeastSignificantZeros().0.leastSignificantOnePosition\ := to_unsigned(0, 16);
                \BitMask::ShiftOutLeastSignificantZeros().0.flag\ := false;
                \BitMask::ShiftOutLeastSignificantZeros().0.return.0\ := to_unsigned(0, 16);
                \BitMask::ShiftOutLeastSignificantZeros().0.binaryOperationResult.0\ := false;
                \BitMask::ShiftOutLeastSignificantZeros().0.binaryOperationResult.1\ := to_signed(0, 32);
            else 
                case \BitMask::ShiftOutLeastSignificantZeros().0._State\ is 
                    when \BitMask::ShiftOutLeastSignificantZeros().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\BitMask::ShiftOutLeastSignificantZeros().0._Started\ = true) then 
                            \BitMask::ShiftOutLeastSignificantZeros().0._State\ := \BitMask::ShiftOutLeastSignificantZeros().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::ShiftOutLeastSignificantZeros().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\BitMask::ShiftOutLeastSignificantZeros().0._Started\ = true) then 
                            \BitMask::ShiftOutLeastSignificantZeros().0._Finished\ <= true;
                        else 
                            \BitMask::ShiftOutLeastSignificantZeros().0._Finished\ <= false;
                            \BitMask::ShiftOutLeastSignificantZeros().0._State\ := \BitMask::ShiftOutLeastSignificantZeros().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::ShiftOutLeastSignificantZeros().0._State_2\ => 
                        \BitMask::ShiftOutLeastSignificantZeros().0.this\ := \BitMask::ShiftOutLeastSignificantZeros().0.this.parameter.In\;
                        -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.BitMask::GetLeastSignificantOnePosition()
                        \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::GetLeastSignificantOnePosition().this.parameter.Out.0\ <= \BitMask::ShiftOutLeastSignificantZeros().0.this\;
                        \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::GetLeastSignificantOnePosition()._Started.0\ <= true;
                        \BitMask::ShiftOutLeastSignificantZeros().0._State\ := \BitMask::ShiftOutLeastSignificantZeros().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::ShiftOutLeastSignificantZeros().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.BitMask::GetLeastSignificantOnePosition()
                        if (\BitMask::ShiftOutLeastSignificantZeros().0.BitMask::GetLeastSignificantOnePosition()._Started.0\ = \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::GetLeastSignificantOnePosition()._Finished.0\) then 
                            \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::GetLeastSignificantOnePosition()._Started.0\ <= false;
                            \BitMask::ShiftOutLeastSignificantZeros().0.return.0\ := \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::GetLeastSignificantOnePosition().return.0\;
                            \BitMask::ShiftOutLeastSignificantZeros().0.leastSignificantOnePosition\ := \BitMask::ShiftOutLeastSignificantZeros().0.return.0\;
                            -- Initializing record fields to their defaults.
                            \BitMask::ShiftOutLeastSignificantZeros().0.bitMask\.\IsNull\ := false;
                            \BitMask::ShiftOutLeastSignificantZeros().0.bitMask\.\Size\ := to_unsigned(0, 16);
                            \BitMask::ShiftOutLeastSignificantZeros().0.bitMask\.\SegmentCount\ := to_unsigned(0, 16);
                            \BitMask::ShiftOutLeastSignificantZeros().0.bitMask\.\Segments\ := (others => to_unsigned(0, 32));
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(Lombiq.Unum.BitMask)
                            \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask).this.parameter.Out.0\ <= \BitMask::ShiftOutLeastSignificantZeros().0.bitMask\;
                            \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask).source.parameter.Out.0\ <= \BitMask::ShiftOutLeastSignificantZeros().0.this\;
                            \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask)._Started.0\ <= true;
                            \BitMask::ShiftOutLeastSignificantZeros().0._State\ := \BitMask::ShiftOutLeastSignificantZeros().0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::ShiftOutLeastSignificantZeros().0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(Lombiq.Unum.BitMask)
                        if (\BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask)._Started.0\ = \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask)._Finished.0\) then 
                            \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask)._Started.0\ <= false;
                            \BitMask::ShiftOutLeastSignificantZeros().0.bitMask\ := \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask).this.parameter.In.0\;
                            \BitMask::ShiftOutLeastSignificantZeros().0.this\ := \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask).source.parameter.In.0\;
                            \BitMask::ShiftOutLeastSignificantZeros().0.binaryOperationResult.0\ := \BitMask::ShiftOutLeastSignificantZeros().0.leastSignificantOnePosition\ = to_unsigned(0, 16);
                            \BitMask::ShiftOutLeastSignificantZeros().0.flag\ := \BitMask::ShiftOutLeastSignificantZeros().0.binaryOperationResult.0\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \BitMask::ShiftOutLeastSignificantZeros().0._State_6\ and ends in state \BitMask::ShiftOutLeastSignificantZeros().0._State_6\.
                            --     * The false branch starts in state \BitMask::ShiftOutLeastSignificantZeros().0._State_7\ and ends in state \BitMask::ShiftOutLeastSignificantZeros().0._State_8\.
                            --     * Execution after either branch will continue in the following state: \BitMask::ShiftOutLeastSignificantZeros().0._State_5\.

                            if (\BitMask::ShiftOutLeastSignificantZeros().0.flag\) then 
                                \BitMask::ShiftOutLeastSignificantZeros().0._State\ := \BitMask::ShiftOutLeastSignificantZeros().0._State_6\;
                            else 
                                \BitMask::ShiftOutLeastSignificantZeros().0._State\ := \BitMask::ShiftOutLeastSignificantZeros().0._State_7\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::ShiftOutLeastSignificantZeros().0._State_5\ => 
                        -- State after the if-else which was started in state \BitMask::ShiftOutLeastSignificantZeros().0._State_4\.
                        \BitMask::ShiftOutLeastSignificantZeros().0.return\ <= \BitMask::ShiftOutLeastSignificantZeros().0.result\;
                        \BitMask::ShiftOutLeastSignificantZeros().0._State\ := \BitMask::ShiftOutLeastSignificantZeros().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::ShiftOutLeastSignificantZeros().0._State_6\ => 
                        -- True branch of the if-else started in state \BitMask::ShiftOutLeastSignificantZeros().0._State_4\.
                        \BitMask::ShiftOutLeastSignificantZeros().0.result\ := \BitMask::ShiftOutLeastSignificantZeros().0.bitMask\;
                        -- Going to the state after the if-else which was started in state \BitMask::ShiftOutLeastSignificantZeros().0._State_4\.
                        if (\BitMask::ShiftOutLeastSignificantZeros().0._State\ = \BitMask::ShiftOutLeastSignificantZeros().0._State_6\) then 
                            \BitMask::ShiftOutLeastSignificantZeros().0._State\ := \BitMask::ShiftOutLeastSignificantZeros().0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::ShiftOutLeastSignificantZeros().0._State_7\ => 
                        -- False branch of the if-else started in state \BitMask::ShiftOutLeastSignificantZeros().0._State_4\.
                        \BitMask::ShiftOutLeastSignificantZeros().0.binaryOperationResult.1\ := resize(signed(\BitMask::ShiftOutLeastSignificantZeros().0.leastSignificantOnePosition\ - to_unsigned(1, 16)), 32);
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_RightShift(Lombiq.Unum.BitMask,System.Int32)
                        \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::op_RightShift(BitMask,Int32).left.parameter.Out.0\ <= \BitMask::ShiftOutLeastSignificantZeros().0.bitMask\;
                        \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::op_RightShift(BitMask,Int32).right.parameter.Out.0\ <= (\BitMask::ShiftOutLeastSignificantZeros().0.binaryOperationResult.1\);
                        \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ <= true;
                        \BitMask::ShiftOutLeastSignificantZeros().0._State\ := \BitMask::ShiftOutLeastSignificantZeros().0._State_8\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::ShiftOutLeastSignificantZeros().0._State_8\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_RightShift(Lombiq.Unum.BitMask,System.Int32)
                        if (\BitMask::ShiftOutLeastSignificantZeros().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ = \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\) then 
                            \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ <= false;
                            \BitMask::ShiftOutLeastSignificantZeros().0.return.1\ := \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::op_RightShift(BitMask,Int32).return.0\;
                            \BitMask::ShiftOutLeastSignificantZeros().0.result\ := \BitMask::ShiftOutLeastSignificantZeros().0.return.1\;
                            -- Going to the state after the if-else which was started in state \BitMask::ShiftOutLeastSignificantZeros().0._State_4\.
                            if (\BitMask::ShiftOutLeastSignificantZeros().0._State\ = \BitMask::ShiftOutLeastSignificantZeros().0._State_8\) then 
                                \BitMask::ShiftOutLeastSignificantZeros().0._State\ := \BitMask::ShiftOutLeastSignificantZeros().0._State_5\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::ShiftOutLeastSignificantZeros().0 state machine end


    -- System.Boolean Lombiq.Unum.BitMask::op_Equality(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 state machine start
    \BitMask::op_Equality(BitMask,BitMask).0._StateMachine\: process (\Clock\) 
        Variable \BitMask::op_Equality(BitMask,BitMask).0._State\: \BitMask::op_Equality(BitMask,BitMask).0._States\ := \BitMask::op_Equality(BitMask,BitMask).0._State_0\;
        Variable \BitMask::op_Equality(BitMask,BitMask).0.left\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_Equality(BitMask,BitMask).0.right\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_Equality(BitMask,BitMask).0.flag\: boolean := false;
        Variable \BitMask::op_Equality(BitMask,BitMask).0.result\: boolean := false;
        Variable \BitMask::op_Equality(BitMask,BitMask).0.num\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_Equality(BitMask,BitMask).0.flag2\: boolean := false;
        Variable \BitMask::op_Equality(BitMask,BitMask).0.binaryOperationResult.0\: boolean := false;
        Variable \BitMask::op_Equality(BitMask,BitMask).0.binaryOperationResult.1\: boolean := false;
        Variable \BitMask::op_Equality(BitMask,BitMask).0.binaryOperationResult.2\: boolean := false;
        Variable \BitMask::op_Equality(BitMask,BitMask).0.binaryOperationResult.3\: boolean := false;
        Variable \BitMask::op_Equality(BitMask,BitMask).0.binaryOperationResult.4\: unsigned(15 downto 0) := to_unsigned(0, 16);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \BitMask::op_Equality(BitMask,BitMask).0._Finished\ <= false;
                \BitMask::op_Equality(BitMask,BitMask).0.return\ <= false;
                \BitMask::op_Equality(BitMask,BitMask).0._State\ := \BitMask::op_Equality(BitMask,BitMask).0._State_0\;
                \BitMask::op_Equality(BitMask,BitMask).0.flag\ := false;
                \BitMask::op_Equality(BitMask,BitMask).0.result\ := false;
                \BitMask::op_Equality(BitMask,BitMask).0.num\ := to_unsigned(0, 16);
                \BitMask::op_Equality(BitMask,BitMask).0.flag2\ := false;
                \BitMask::op_Equality(BitMask,BitMask).0.binaryOperationResult.0\ := false;
                \BitMask::op_Equality(BitMask,BitMask).0.binaryOperationResult.1\ := false;
                \BitMask::op_Equality(BitMask,BitMask).0.binaryOperationResult.2\ := false;
                \BitMask::op_Equality(BitMask,BitMask).0.binaryOperationResult.3\ := false;
                \BitMask::op_Equality(BitMask,BitMask).0.binaryOperationResult.4\ := to_unsigned(0, 16);
            else 
                case \BitMask::op_Equality(BitMask,BitMask).0._State\ is 
                    when \BitMask::op_Equality(BitMask,BitMask).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\BitMask::op_Equality(BitMask,BitMask).0._Started\ = true) then 
                            \BitMask::op_Equality(BitMask,BitMask).0._State\ := \BitMask::op_Equality(BitMask,BitMask).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Equality(BitMask,BitMask).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\BitMask::op_Equality(BitMask,BitMask).0._Started\ = true) then 
                            \BitMask::op_Equality(BitMask,BitMask).0._Finished\ <= true;
                        else 
                            \BitMask::op_Equality(BitMask,BitMask).0._Finished\ <= false;
                            \BitMask::op_Equality(BitMask,BitMask).0._State\ := \BitMask::op_Equality(BitMask,BitMask).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Equality(BitMask,BitMask).0._State_2\ => 
                        \BitMask::op_Equality(BitMask,BitMask).0.left\ := \BitMask::op_Equality(BitMask,BitMask).0.left.parameter.In\;
                        \BitMask::op_Equality(BitMask,BitMask).0.right\ := \BitMask::op_Equality(BitMask,BitMask).0.right.parameter.In\;
                        \BitMask::op_Equality(BitMask,BitMask).0.binaryOperationResult.0\ := \BitMask::op_Equality(BitMask,BitMask).0.left\.\SegmentCount\ /= \BitMask::op_Equality(BitMask,BitMask).0.right\.\SegmentCount\;
                        \BitMask::op_Equality(BitMask,BitMask).0.flag\ := \BitMask::op_Equality(BitMask,BitMask).0.binaryOperationResult.0\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::op_Equality(BitMask,BitMask).0._State_4\ and ends in state \BitMask::op_Equality(BitMask,BitMask).0._State_4\.
                        --     * The false branch starts in state \BitMask::op_Equality(BitMask,BitMask).0._State_5\ and ends in state \BitMask::op_Equality(BitMask,BitMask).0._State_7\.
                        --     * Execution after either branch will continue in the following state: \BitMask::op_Equality(BitMask,BitMask).0._State_3\.

                        if (\BitMask::op_Equality(BitMask,BitMask).0.flag\) then 
                            \BitMask::op_Equality(BitMask,BitMask).0._State\ := \BitMask::op_Equality(BitMask,BitMask).0._State_4\;
                        else 
                            \BitMask::op_Equality(BitMask,BitMask).0._State\ := \BitMask::op_Equality(BitMask,BitMask).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_Equality(BitMask,BitMask).0._State_3\ => 
                        -- State after the if-else which was started in state \BitMask::op_Equality(BitMask,BitMask).0._State_2\.
                        \BitMask::op_Equality(BitMask,BitMask).0.return\ <= \BitMask::op_Equality(BitMask,BitMask).0.result\;
                        \BitMask::op_Equality(BitMask,BitMask).0._State\ := \BitMask::op_Equality(BitMask,BitMask).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Equality(BitMask,BitMask).0._State_4\ => 
                        -- True branch of the if-else started in state \BitMask::op_Equality(BitMask,BitMask).0._State_2\.
                        \BitMask::op_Equality(BitMask,BitMask).0.result\ := False;
                        -- Going to the state after the if-else which was started in state \BitMask::op_Equality(BitMask,BitMask).0._State_2\.
                        if (\BitMask::op_Equality(BitMask,BitMask).0._State\ = \BitMask::op_Equality(BitMask,BitMask).0._State_4\) then 
                            \BitMask::op_Equality(BitMask,BitMask).0._State\ := \BitMask::op_Equality(BitMask,BitMask).0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Equality(BitMask,BitMask).0._State_5\ => 
                        -- False branch of the if-else started in state \BitMask::op_Equality(BitMask,BitMask).0._State_2\.
                        \BitMask::op_Equality(BitMask,BitMask).0.num\ := to_unsigned(0, 16);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \BitMask::op_Equality(BitMask,BitMask).0.binaryOperationResult.1\ := \BitMask::op_Equality(BitMask,BitMask).0.num\ < \BitMask::op_Equality(BitMask,BitMask).0.left\.\SegmentCount\;
                        if (\BitMask::op_Equality(BitMask,BitMask).0.binaryOperationResult.1\) then 
                            \BitMask::op_Equality(BitMask,BitMask).0._State\ := \BitMask::op_Equality(BitMask,BitMask).0._State_6\;
                        else 
                            \BitMask::op_Equality(BitMask,BitMask).0._State\ := \BitMask::op_Equality(BitMask,BitMask).0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_Equality(BitMask,BitMask).0._State_6\ => 
                        -- Repeated state of the while loop which was started in state \BitMask::op_Equality(BitMask,BitMask).0._State_5\.
                        -- The while loop's condition:
                        \BitMask::op_Equality(BitMask,BitMask).0.binaryOperationResult.2\ := \BitMask::op_Equality(BitMask,BitMask).0.num\ < \BitMask::op_Equality(BitMask,BitMask).0.left\.\SegmentCount\;
                        if (\BitMask::op_Equality(BitMask,BitMask).0.binaryOperationResult.2\) then 
                            \BitMask::op_Equality(BitMask,BitMask).0.binaryOperationResult.3\ := \BitMask::op_Equality(BitMask,BitMask).0.left\.\Segments\(to_integer(resize(signed(\BitMask::op_Equality(BitMask,BitMask).0.num\), 32))) /= \BitMask::op_Equality(BitMask,BitMask).0.right\.\Segments\(to_integer(resize(signed(\BitMask::op_Equality(BitMask,BitMask).0.num\), 32)));
                            \BitMask::op_Equality(BitMask,BitMask).0.flag2\ := \BitMask::op_Equality(BitMask,BitMask).0.binaryOperationResult.3\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \BitMask::op_Equality(BitMask,BitMask).0._State_9\ and ends in state \BitMask::op_Equality(BitMask,BitMask).0._State_9\.
                            --     * Execution after either branch will continue in the following state: \BitMask::op_Equality(BitMask,BitMask).0._State_8\.

                            if (\BitMask::op_Equality(BitMask,BitMask).0.flag2\) then 
                                \BitMask::op_Equality(BitMask,BitMask).0._State\ := \BitMask::op_Equality(BitMask,BitMask).0._State_9\;
                            else 
                                -- There was no false branch, so going directly to the state after the if-else.
                                \BitMask::op_Equality(BitMask,BitMask).0._State\ := \BitMask::op_Equality(BitMask,BitMask).0._State_8\;
                            end if;
                        else 
                            \BitMask::op_Equality(BitMask,BitMask).0._State\ := \BitMask::op_Equality(BitMask,BitMask).0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \BitMask::op_Equality(BitMask,BitMask).0._State_7\ => 
                        -- State after the while loop which was started in state \BitMask::op_Equality(BitMask,BitMask).0._State_5\.
                        \BitMask::op_Equality(BitMask,BitMask).0.result\ := True;
                        -- Going to the state after the if-else which was started in state \BitMask::op_Equality(BitMask,BitMask).0._State_2\.
                        if (\BitMask::op_Equality(BitMask,BitMask).0._State\ = \BitMask::op_Equality(BitMask,BitMask).0._State_7\) then 
                            \BitMask::op_Equality(BitMask,BitMask).0._State\ := \BitMask::op_Equality(BitMask,BitMask).0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Equality(BitMask,BitMask).0._State_8\ => 
                        -- State after the if-else which was started in state \BitMask::op_Equality(BitMask,BitMask).0._State_6\.
                        \BitMask::op_Equality(BitMask,BitMask).0.binaryOperationResult.4\ := \BitMask::op_Equality(BitMask,BitMask).0.num\ + to_unsigned(1, 16);
                        \BitMask::op_Equality(BitMask,BitMask).0.num\ := \BitMask::op_Equality(BitMask,BitMask).0.binaryOperationResult.4\;
                        -- Returning to the repeated state of the while loop which was started in state \BitMask::op_Equality(BitMask,BitMask).0._State_5\ if the loop wasn't exited with a state change.
                        if (\BitMask::op_Equality(BitMask,BitMask).0._State\ = \BitMask::op_Equality(BitMask,BitMask).0._State_8\) then 
                            \BitMask::op_Equality(BitMask,BitMask).0._State\ := \BitMask::op_Equality(BitMask,BitMask).0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_Equality(BitMask,BitMask).0._State_9\ => 
                        -- True branch of the if-else started in state \BitMask::op_Equality(BitMask,BitMask).0._State_6\.
                        \BitMask::op_Equality(BitMask,BitMask).0.result\ := False;
                        \BitMask::op_Equality(BitMask,BitMask).0.return\ <= \BitMask::op_Equality(BitMask,BitMask).0.result\;
                        \BitMask::op_Equality(BitMask,BitMask).0._State\ := \BitMask::op_Equality(BitMask,BitMask).0._State_1\;
                        -- Going to the state after the if-else which was started in state \BitMask::op_Equality(BitMask,BitMask).0._State_6\.
                        if (\BitMask::op_Equality(BitMask,BitMask).0._State\ = \BitMask::op_Equality(BitMask,BitMask).0._State_9\) then 
                            \BitMask::op_Equality(BitMask,BitMask).0._State\ := \BitMask::op_Equality(BitMask,BitMask).0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Lombiq.Unum.BitMask::op_Equality(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 state machine end


    -- System.Boolean Lombiq.Unum.BitMask::op_GreaterThan(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 state machine start
    \BitMask::op_GreaterThan(BitMask,BitMask).0._StateMachine\: process (\Clock\) 
        Variable \BitMask::op_GreaterThan(BitMask,BitMask).0._State\: \BitMask::op_GreaterThan(BitMask,BitMask).0._States\ := \BitMask::op_GreaterThan(BitMask,BitMask).0._State_0\;
        Variable \BitMask::op_GreaterThan(BitMask,BitMask).0.left\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_GreaterThan(BitMask,BitMask).0.right\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_GreaterThan(BitMask,BitMask).0.num\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_GreaterThan(BitMask,BitMask).0.flag\: boolean := false;
        Variable \BitMask::op_GreaterThan(BitMask,BitMask).0.result\: boolean := false;
        Variable \BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.0\: boolean := false;
        Variable \BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.1\: boolean := false;
        Variable \BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.3\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.4\: boolean := false;
        Variable \BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.5\: unsigned(15 downto 0) := to_unsigned(0, 16);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \BitMask::op_GreaterThan(BitMask,BitMask).0._Finished\ <= false;
                \BitMask::op_GreaterThan(BitMask,BitMask).0.return\ <= false;
                \BitMask::op_GreaterThan(BitMask,BitMask).0._State\ := \BitMask::op_GreaterThan(BitMask,BitMask).0._State_0\;
                \BitMask::op_GreaterThan(BitMask,BitMask).0.num\ := to_unsigned(0, 16);
                \BitMask::op_GreaterThan(BitMask,BitMask).0.flag\ := false;
                \BitMask::op_GreaterThan(BitMask,BitMask).0.result\ := false;
                \BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.0\ := false;
                \BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.1\ := false;
                \BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.2\ := to_signed(0, 32);
                \BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.3\ := to_signed(0, 32);
                \BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.4\ := false;
                \BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.5\ := to_unsigned(0, 16);
            else 
                case \BitMask::op_GreaterThan(BitMask,BitMask).0._State\ is 
                    when \BitMask::op_GreaterThan(BitMask,BitMask).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\BitMask::op_GreaterThan(BitMask,BitMask).0._Started\ = true) then 
                            \BitMask::op_GreaterThan(BitMask,BitMask).0._State\ := \BitMask::op_GreaterThan(BitMask,BitMask).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_GreaterThan(BitMask,BitMask).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\BitMask::op_GreaterThan(BitMask,BitMask).0._Started\ = true) then 
                            \BitMask::op_GreaterThan(BitMask,BitMask).0._Finished\ <= true;
                        else 
                            \BitMask::op_GreaterThan(BitMask,BitMask).0._Finished\ <= false;
                            \BitMask::op_GreaterThan(BitMask,BitMask).0._State\ := \BitMask::op_GreaterThan(BitMask,BitMask).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_GreaterThan(BitMask,BitMask).0._State_2\ => 
                        \BitMask::op_GreaterThan(BitMask,BitMask).0.left\ := \BitMask::op_GreaterThan(BitMask,BitMask).0.left.parameter.In\;
                        \BitMask::op_GreaterThan(BitMask,BitMask).0.right\ := \BitMask::op_GreaterThan(BitMask,BitMask).0.right.parameter.In\;
                        \BitMask::op_GreaterThan(BitMask,BitMask).0.num\ := to_unsigned(1, 16);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.0\ := \BitMask::op_GreaterThan(BitMask,BitMask).0.num\ <= \BitMask::op_GreaterThan(BitMask,BitMask).0.left\.\SegmentCount\;
                        if (\BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.0\) then 
                            \BitMask::op_GreaterThan(BitMask,BitMask).0._State\ := \BitMask::op_GreaterThan(BitMask,BitMask).0._State_3\;
                        else 
                            \BitMask::op_GreaterThan(BitMask,BitMask).0._State\ := \BitMask::op_GreaterThan(BitMask,BitMask).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_GreaterThan(BitMask,BitMask).0._State_3\ => 
                        -- Repeated state of the while loop which was started in state \BitMask::op_GreaterThan(BitMask,BitMask).0._State_2\.
                        -- The while loop's condition:
                        \BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.1\ := \BitMask::op_GreaterThan(BitMask,BitMask).0.num\ <= \BitMask::op_GreaterThan(BitMask,BitMask).0.left\.\SegmentCount\;
                        if (\BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.1\) then 
                            \BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.2\ := resize(signed(\BitMask::op_GreaterThan(BitMask,BitMask).0.left\.\SegmentCount\ - \BitMask::op_GreaterThan(BitMask,BitMask).0.num\), 32);
                            \BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.3\ := resize(signed(\BitMask::op_GreaterThan(BitMask,BitMask).0.left\.\SegmentCount\ - \BitMask::op_GreaterThan(BitMask,BitMask).0.num\), 32);
                            \BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.4\ := \BitMask::op_GreaterThan(BitMask,BitMask).0.left\.\Segments\(to_integer((\BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.2\))) > \BitMask::op_GreaterThan(BitMask,BitMask).0.right\.\Segments\(to_integer((\BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.3\)));
                            \BitMask::op_GreaterThan(BitMask,BitMask).0.flag\ := \BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.4\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \BitMask::op_GreaterThan(BitMask,BitMask).0._State_6\ and ends in state \BitMask::op_GreaterThan(BitMask,BitMask).0._State_6\.
                            --     * Execution after either branch will continue in the following state: \BitMask::op_GreaterThan(BitMask,BitMask).0._State_5\.

                            if (\BitMask::op_GreaterThan(BitMask,BitMask).0.flag\) then 
                                \BitMask::op_GreaterThan(BitMask,BitMask).0._State\ := \BitMask::op_GreaterThan(BitMask,BitMask).0._State_6\;
                            else 
                                -- There was no false branch, so going directly to the state after the if-else.
                                \BitMask::op_GreaterThan(BitMask,BitMask).0._State\ := \BitMask::op_GreaterThan(BitMask,BitMask).0._State_5\;
                            end if;
                        else 
                            \BitMask::op_GreaterThan(BitMask,BitMask).0._State\ := \BitMask::op_GreaterThan(BitMask,BitMask).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.4
                    when \BitMask::op_GreaterThan(BitMask,BitMask).0._State_4\ => 
                        -- State after the while loop which was started in state \BitMask::op_GreaterThan(BitMask,BitMask).0._State_2\.
                        \BitMask::op_GreaterThan(BitMask,BitMask).0.result\ := False;
                        \BitMask::op_GreaterThan(BitMask,BitMask).0.return\ <= False;
                        \BitMask::op_GreaterThan(BitMask,BitMask).0._State\ := \BitMask::op_GreaterThan(BitMask,BitMask).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_GreaterThan(BitMask,BitMask).0._State_5\ => 
                        -- State after the if-else which was started in state \BitMask::op_GreaterThan(BitMask,BitMask).0._State_3\.
                        \BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.5\ := \BitMask::op_GreaterThan(BitMask,BitMask).0.num\ + to_unsigned(1, 16);
                        \BitMask::op_GreaterThan(BitMask,BitMask).0.num\ := \BitMask::op_GreaterThan(BitMask,BitMask).0.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \BitMask::op_GreaterThan(BitMask,BitMask).0._State_2\ if the loop wasn't exited with a state change.
                        if (\BitMask::op_GreaterThan(BitMask,BitMask).0._State\ = \BitMask::op_GreaterThan(BitMask,BitMask).0._State_5\) then 
                            \BitMask::op_GreaterThan(BitMask,BitMask).0._State\ := \BitMask::op_GreaterThan(BitMask,BitMask).0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_GreaterThan(BitMask,BitMask).0._State_6\ => 
                        -- True branch of the if-else started in state \BitMask::op_GreaterThan(BitMask,BitMask).0._State_3\.
                        \BitMask::op_GreaterThan(BitMask,BitMask).0.result\ := True;
                        \BitMask::op_GreaterThan(BitMask,BitMask).0.return\ <= \BitMask::op_GreaterThan(BitMask,BitMask).0.result\;
                        \BitMask::op_GreaterThan(BitMask,BitMask).0._State\ := \BitMask::op_GreaterThan(BitMask,BitMask).0._State_1\;
                        -- Going to the state after the if-else which was started in state \BitMask::op_GreaterThan(BitMask,BitMask).0._State_3\.
                        if (\BitMask::op_GreaterThan(BitMask,BitMask).0._State\ = \BitMask::op_GreaterThan(BitMask,BitMask).0._State_6\) then 
                            \BitMask::op_GreaterThan(BitMask,BitMask).0._State\ := \BitMask::op_GreaterThan(BitMask,BitMask).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Lombiq.Unum.BitMask::op_GreaterThan(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 state machine end


    -- System.Boolean Lombiq.Unum.BitMask::op_LessThan(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 state machine start
    \BitMask::op_LessThan(BitMask,BitMask).0._StateMachine\: process (\Clock\) 
        Variable \BitMask::op_LessThan(BitMask,BitMask).0._State\: \BitMask::op_LessThan(BitMask,BitMask).0._States\ := \BitMask::op_LessThan(BitMask,BitMask).0._State_0\;
        Variable \BitMask::op_LessThan(BitMask,BitMask).0.left\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_LessThan(BitMask,BitMask).0.right\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_LessThan(BitMask,BitMask).0.num\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_LessThan(BitMask,BitMask).0.flag\: boolean := false;
        Variable \BitMask::op_LessThan(BitMask,BitMask).0.result\: boolean := false;
        Variable \BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.0\: boolean := false;
        Variable \BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.1\: boolean := false;
        Variable \BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.3\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.4\: boolean := false;
        Variable \BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.5\: unsigned(15 downto 0) := to_unsigned(0, 16);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \BitMask::op_LessThan(BitMask,BitMask).0._Finished\ <= false;
                \BitMask::op_LessThan(BitMask,BitMask).0.return\ <= false;
                \BitMask::op_LessThan(BitMask,BitMask).0._State\ := \BitMask::op_LessThan(BitMask,BitMask).0._State_0\;
                \BitMask::op_LessThan(BitMask,BitMask).0.num\ := to_unsigned(0, 16);
                \BitMask::op_LessThan(BitMask,BitMask).0.flag\ := false;
                \BitMask::op_LessThan(BitMask,BitMask).0.result\ := false;
                \BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.0\ := false;
                \BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.1\ := false;
                \BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.2\ := to_signed(0, 32);
                \BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.3\ := to_signed(0, 32);
                \BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.4\ := false;
                \BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.5\ := to_unsigned(0, 16);
            else 
                case \BitMask::op_LessThan(BitMask,BitMask).0._State\ is 
                    when \BitMask::op_LessThan(BitMask,BitMask).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\BitMask::op_LessThan(BitMask,BitMask).0._Started\ = true) then 
                            \BitMask::op_LessThan(BitMask,BitMask).0._State\ := \BitMask::op_LessThan(BitMask,BitMask).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_LessThan(BitMask,BitMask).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\BitMask::op_LessThan(BitMask,BitMask).0._Started\ = true) then 
                            \BitMask::op_LessThan(BitMask,BitMask).0._Finished\ <= true;
                        else 
                            \BitMask::op_LessThan(BitMask,BitMask).0._Finished\ <= false;
                            \BitMask::op_LessThan(BitMask,BitMask).0._State\ := \BitMask::op_LessThan(BitMask,BitMask).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_LessThan(BitMask,BitMask).0._State_2\ => 
                        \BitMask::op_LessThan(BitMask,BitMask).0.left\ := \BitMask::op_LessThan(BitMask,BitMask).0.left.parameter.In\;
                        \BitMask::op_LessThan(BitMask,BitMask).0.right\ := \BitMask::op_LessThan(BitMask,BitMask).0.right.parameter.In\;
                        \BitMask::op_LessThan(BitMask,BitMask).0.num\ := to_unsigned(1, 16);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.0\ := \BitMask::op_LessThan(BitMask,BitMask).0.num\ <= \BitMask::op_LessThan(BitMask,BitMask).0.left\.\SegmentCount\;
                        if (\BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.0\) then 
                            \BitMask::op_LessThan(BitMask,BitMask).0._State\ := \BitMask::op_LessThan(BitMask,BitMask).0._State_3\;
                        else 
                            \BitMask::op_LessThan(BitMask,BitMask).0._State\ := \BitMask::op_LessThan(BitMask,BitMask).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_LessThan(BitMask,BitMask).0._State_3\ => 
                        -- Repeated state of the while loop which was started in state \BitMask::op_LessThan(BitMask,BitMask).0._State_2\.
                        -- The while loop's condition:
                        \BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.1\ := \BitMask::op_LessThan(BitMask,BitMask).0.num\ <= \BitMask::op_LessThan(BitMask,BitMask).0.left\.\SegmentCount\;
                        if (\BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.1\) then 
                            \BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.2\ := resize(signed(\BitMask::op_LessThan(BitMask,BitMask).0.left\.\SegmentCount\ - \BitMask::op_LessThan(BitMask,BitMask).0.num\), 32);
                            \BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.3\ := resize(signed(\BitMask::op_LessThan(BitMask,BitMask).0.left\.\SegmentCount\ - \BitMask::op_LessThan(BitMask,BitMask).0.num\), 32);
                            \BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.4\ := \BitMask::op_LessThan(BitMask,BitMask).0.left\.\Segments\(to_integer((\BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.2\))) < \BitMask::op_LessThan(BitMask,BitMask).0.right\.\Segments\(to_integer((\BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.3\)));
                            \BitMask::op_LessThan(BitMask,BitMask).0.flag\ := \BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.4\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \BitMask::op_LessThan(BitMask,BitMask).0._State_6\ and ends in state \BitMask::op_LessThan(BitMask,BitMask).0._State_6\.
                            --     * Execution after either branch will continue in the following state: \BitMask::op_LessThan(BitMask,BitMask).0._State_5\.

                            if (\BitMask::op_LessThan(BitMask,BitMask).0.flag\) then 
                                \BitMask::op_LessThan(BitMask,BitMask).0._State\ := \BitMask::op_LessThan(BitMask,BitMask).0._State_6\;
                            else 
                                -- There was no false branch, so going directly to the state after the if-else.
                                \BitMask::op_LessThan(BitMask,BitMask).0._State\ := \BitMask::op_LessThan(BitMask,BitMask).0._State_5\;
                            end if;
                        else 
                            \BitMask::op_LessThan(BitMask,BitMask).0._State\ := \BitMask::op_LessThan(BitMask,BitMask).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.4
                    when \BitMask::op_LessThan(BitMask,BitMask).0._State_4\ => 
                        -- State after the while loop which was started in state \BitMask::op_LessThan(BitMask,BitMask).0._State_2\.
                        \BitMask::op_LessThan(BitMask,BitMask).0.result\ := False;
                        \BitMask::op_LessThan(BitMask,BitMask).0.return\ <= False;
                        \BitMask::op_LessThan(BitMask,BitMask).0._State\ := \BitMask::op_LessThan(BitMask,BitMask).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_LessThan(BitMask,BitMask).0._State_5\ => 
                        -- State after the if-else which was started in state \BitMask::op_LessThan(BitMask,BitMask).0._State_3\.
                        \BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.5\ := \BitMask::op_LessThan(BitMask,BitMask).0.num\ + to_unsigned(1, 16);
                        \BitMask::op_LessThan(BitMask,BitMask).0.num\ := \BitMask::op_LessThan(BitMask,BitMask).0.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \BitMask::op_LessThan(BitMask,BitMask).0._State_2\ if the loop wasn't exited with a state change.
                        if (\BitMask::op_LessThan(BitMask,BitMask).0._State\ = \BitMask::op_LessThan(BitMask,BitMask).0._State_5\) then 
                            \BitMask::op_LessThan(BitMask,BitMask).0._State\ := \BitMask::op_LessThan(BitMask,BitMask).0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_LessThan(BitMask,BitMask).0._State_6\ => 
                        -- True branch of the if-else started in state \BitMask::op_LessThan(BitMask,BitMask).0._State_3\.
                        \BitMask::op_LessThan(BitMask,BitMask).0.result\ := True;
                        \BitMask::op_LessThan(BitMask,BitMask).0.return\ <= \BitMask::op_LessThan(BitMask,BitMask).0.result\;
                        \BitMask::op_LessThan(BitMask,BitMask).0._State\ := \BitMask::op_LessThan(BitMask,BitMask).0._State_1\;
                        -- Going to the state after the if-else which was started in state \BitMask::op_LessThan(BitMask,BitMask).0._State_3\.
                        if (\BitMask::op_LessThan(BitMask,BitMask).0._State\ = \BitMask::op_LessThan(BitMask,BitMask).0._State_6\) then 
                            \BitMask::op_LessThan(BitMask,BitMask).0._State\ := \BitMask::op_LessThan(BitMask,BitMask).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Lombiq.Unum.BitMask::op_LessThan(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 state machine end


    -- System.Boolean Lombiq.Unum.BitMask::op_GreaterThanOrEqual(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 state machine start
    \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._StateMachine\: process (\Clock\) 
        Variable \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._State\: \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._States\ := \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._State_0\;
        Variable \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.left\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.right\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.return.0\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._Finished\ <= false;
                \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.return\ <= false;
                \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.BitMask::op_LessThan(BitMask,BitMask)._Started.0\ <= false;
                \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._State\ := \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._State_0\;
                \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.return.0\ := false;
            else 
                case \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._State\ is 
                    when \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._Started\ = true) then 
                            \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._State\ := \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._Started\ = true) then 
                            \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._Finished\ <= true;
                        else 
                            \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._Finished\ <= false;
                            \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._State\ := \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._State_2\ => 
                        \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.left\ := \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.left.parameter.In\;
                        \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.right\ := \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.right.parameter.In\;
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.BitMask::op_LessThan(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.BitMask::op_LessThan(BitMask,BitMask).left.parameter.Out.0\ <= \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.left\;
                        \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.BitMask::op_LessThan(BitMask,BitMask).right.parameter.Out.0\ <= \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.right\;
                        \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.BitMask::op_LessThan(BitMask,BitMask)._Started.0\ <= true;
                        \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._State\ := \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.BitMask::op_LessThan(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.BitMask::op_LessThan(BitMask,BitMask)._Started.0\ = \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.BitMask::op_LessThan(BitMask,BitMask)._Finished.0\) then 
                            \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.BitMask::op_LessThan(BitMask,BitMask)._Started.0\ <= false;
                            \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.return.0\ := \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.BitMask::op_LessThan(BitMask,BitMask).return.0\;
                            \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.return\ <= not(\BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.return.0\);
                            \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._State\ := \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Lombiq.Unum.BitMask::op_GreaterThanOrEqual(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,System.UInt32).0 state machine start
    \BitMask::op_Addition(BitMask,UInt32).0._StateMachine\: process (\Clock\) 
        Variable \BitMask::op_Addition(BitMask,UInt32).0._State\: \BitMask::op_Addition(BitMask,UInt32).0._States\ := \BitMask::op_Addition(BitMask,UInt32).0._State_0\;
        Variable \BitMask::op_Addition(BitMask,UInt32).0.left\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_Addition(BitMask,UInt32).0.right\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_Addition(BitMask,UInt32).0.array354f1c9f95760fbd3aea950ed967f55dcf8694b14f050cae5da73e6d4fbc0271\: \unsigned32_Array\(0 to 0) := (others => to_unsigned(0, 32));
        Variable \BitMask::op_Addition(BitMask,UInt32).0.object318df7b6a8d78dabf5d944006517b7f614152baa1ab93d6683e48e42bf520fd3\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_Addition(BitMask,UInt32).0.return.0\: \Lombiq.Unum.BitMask\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \BitMask::op_Addition(BitMask,UInt32).0._Finished\ <= false;
                \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 32));
                \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                \BitMask::op_Addition(BitMask,UInt32).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= false;
                \BitMask::op_Addition(BitMask,UInt32).0._State\ := \BitMask::op_Addition(BitMask,UInt32).0._State_0\;
                \BitMask::op_Addition(BitMask,UInt32).0.right\ := to_unsigned(0, 32);
                \BitMask::op_Addition(BitMask,UInt32).0.array354f1c9f95760fbd3aea950ed967f55dcf8694b14f050cae5da73e6d4fbc0271\ := (others => to_unsigned(0, 32));
            else 
                case \BitMask::op_Addition(BitMask,UInt32).0._State\ is 
                    when \BitMask::op_Addition(BitMask,UInt32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\BitMask::op_Addition(BitMask,UInt32).0._Started\ = true) then 
                            \BitMask::op_Addition(BitMask,UInt32).0._State\ := \BitMask::op_Addition(BitMask,UInt32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Addition(BitMask,UInt32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\BitMask::op_Addition(BitMask,UInt32).0._Started\ = true) then 
                            \BitMask::op_Addition(BitMask,UInt32).0._Finished\ <= true;
                        else 
                            \BitMask::op_Addition(BitMask,UInt32).0._Finished\ <= false;
                            \BitMask::op_Addition(BitMask,UInt32).0._State\ := \BitMask::op_Addition(BitMask,UInt32).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Addition(BitMask,UInt32).0._State_2\ => 
                        \BitMask::op_Addition(BitMask,UInt32).0.left\ := \BitMask::op_Addition(BitMask,UInt32).0.left.parameter.In\;
                        \BitMask::op_Addition(BitMask,UInt32).0.right\ := \BitMask::op_Addition(BitMask,UInt32).0.right.parameter.In\;
                        \BitMask::op_Addition(BitMask,UInt32).0.array354f1c9f95760fbd3aea950ed967f55dcf8694b14f050cae5da73e6d4fbc0271\ := (others => to_unsigned(0, 32));
                        \BitMask::op_Addition(BitMask,UInt32).0.array354f1c9f95760fbd3aea950ed967f55dcf8694b14f050cae5da73e6d4fbc0271\(to_integer(to_signed(0, 32))) := \BitMask::op_Addition(BitMask,UInt32).0.right\;
                        -- Initializing record fields to their defaults.
                        \BitMask::op_Addition(BitMask,UInt32).0.object318df7b6a8d78dabf5d944006517b7f614152baa1ab93d6683e48e42bf520fd3\.\IsNull\ := false;
                        \BitMask::op_Addition(BitMask,UInt32).0.object318df7b6a8d78dabf5d944006517b7f614152baa1ab93d6683e48e42bf520fd3\.\Size\ := to_unsigned(0, 16);
                        \BitMask::op_Addition(BitMask,UInt32).0.object318df7b6a8d78dabf5d944006517b7f614152baa1ab93d6683e48e42bf520fd3\.\SegmentCount\ := to_unsigned(0, 16);
                        \BitMask::op_Addition(BitMask,UInt32).0.object318df7b6a8d78dabf5d944006517b7f614152baa1ab93d6683e48e42bf520fd3\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\ <= \BitMask::op_Addition(BitMask,UInt32).0.object318df7b6a8d78dabf5d944006517b7f614152baa1ab93d6683e48e42bf520fd3\;
                        \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\(0 to 0) <= \BitMask::op_Addition(BitMask,UInt32).0.array354f1c9f95760fbd3aea950ed967f55dcf8694b14f050cae5da73e6d4fbc0271\;
                        \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= \BitMask::op_Addition(BitMask,UInt32).0.left\.\Size\;
                        \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= true;
                        \BitMask::op_Addition(BitMask,UInt32).0._State\ := \BitMask::op_Addition(BitMask,UInt32).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Addition(BitMask,UInt32).0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        if (\BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\) then 
                            \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                            \BitMask::op_Addition(BitMask,UInt32).0.object318df7b6a8d78dabf5d944006517b7f614152baa1ab93d6683e48e42bf520fd3\ := \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\;
                            \BitMask::op_Addition(BitMask,UInt32).0.array354f1c9f95760fbd3aea950ed967f55dcf8694b14f050cae5da73e6d4fbc0271\ := \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\(0 to 0);
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \BitMask::op_Addition(BitMask,UInt32).0.BitMask::op_Addition(BitMask,BitMask).left.parameter.Out.0\ <= \BitMask::op_Addition(BitMask,UInt32).0.left\;
                            \BitMask::op_Addition(BitMask,UInt32).0.BitMask::op_Addition(BitMask,BitMask).right.parameter.Out.0\ <= \BitMask::op_Addition(BitMask,UInt32).0.object318df7b6a8d78dabf5d944006517b7f614152baa1ab93d6683e48e42bf520fd3\;
                            \BitMask::op_Addition(BitMask,UInt32).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= true;
                            \BitMask::op_Addition(BitMask,UInt32).0._State\ := \BitMask::op_Addition(BitMask,UInt32).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Addition(BitMask,UInt32).0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\BitMask::op_Addition(BitMask,UInt32).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ = \BitMask::op_Addition(BitMask,UInt32).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\) then 
                            \BitMask::op_Addition(BitMask,UInt32).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= false;
                            \BitMask::op_Addition(BitMask,UInt32).0.return.0\ := \BitMask::op_Addition(BitMask,UInt32).0.BitMask::op_Addition(BitMask,BitMask).return.0\;
                            \BitMask::op_Addition(BitMask,UInt32).0.return\ <= \BitMask::op_Addition(BitMask,UInt32).0.return.0\;
                            \BitMask::op_Addition(BitMask,UInt32).0._State\ := \BitMask::op_Addition(BitMask,UInt32).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,System.UInt32).0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,System.UInt32).0 state machine start
    \BitMask::op_Subtraction(BitMask,UInt32).0._StateMachine\: process (\Clock\) 
        Variable \BitMask::op_Subtraction(BitMask,UInt32).0._State\: \BitMask::op_Subtraction(BitMask,UInt32).0._States\ := \BitMask::op_Subtraction(BitMask,UInt32).0._State_0\;
        Variable \BitMask::op_Subtraction(BitMask,UInt32).0.left\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_Subtraction(BitMask,UInt32).0.right\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_Subtraction(BitMask,UInt32).0.arrayc8aa351a91a705be1462d4711470c40b589d09135c08d50b79a45acfa9e94d27\: \unsigned32_Array\(0 to 0) := (others => to_unsigned(0, 32));
        Variable \BitMask::op_Subtraction(BitMask,UInt32).0.object77d16c4ef26cad24ef177b742166d622e968246a8b3c1e923c73e932760e2cc3\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_Subtraction(BitMask,UInt32).0.return.0\: \Lombiq.Unum.BitMask\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \BitMask::op_Subtraction(BitMask,UInt32).0._Finished\ <= false;
                \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 32));
                \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ <= false;
                \BitMask::op_Subtraction(BitMask,UInt32).0._State\ := \BitMask::op_Subtraction(BitMask,UInt32).0._State_0\;
                \BitMask::op_Subtraction(BitMask,UInt32).0.right\ := to_unsigned(0, 32);
                \BitMask::op_Subtraction(BitMask,UInt32).0.arrayc8aa351a91a705be1462d4711470c40b589d09135c08d50b79a45acfa9e94d27\ := (others => to_unsigned(0, 32));
            else 
                case \BitMask::op_Subtraction(BitMask,UInt32).0._State\ is 
                    when \BitMask::op_Subtraction(BitMask,UInt32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\BitMask::op_Subtraction(BitMask,UInt32).0._Started\ = true) then 
                            \BitMask::op_Subtraction(BitMask,UInt32).0._State\ := \BitMask::op_Subtraction(BitMask,UInt32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Subtraction(BitMask,UInt32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\BitMask::op_Subtraction(BitMask,UInt32).0._Started\ = true) then 
                            \BitMask::op_Subtraction(BitMask,UInt32).0._Finished\ <= true;
                        else 
                            \BitMask::op_Subtraction(BitMask,UInt32).0._Finished\ <= false;
                            \BitMask::op_Subtraction(BitMask,UInt32).0._State\ := \BitMask::op_Subtraction(BitMask,UInt32).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Subtraction(BitMask,UInt32).0._State_2\ => 
                        \BitMask::op_Subtraction(BitMask,UInt32).0.left\ := \BitMask::op_Subtraction(BitMask,UInt32).0.left.parameter.In\;
                        \BitMask::op_Subtraction(BitMask,UInt32).0.right\ := \BitMask::op_Subtraction(BitMask,UInt32).0.right.parameter.In\;
                        \BitMask::op_Subtraction(BitMask,UInt32).0.arrayc8aa351a91a705be1462d4711470c40b589d09135c08d50b79a45acfa9e94d27\ := (others => to_unsigned(0, 32));
                        \BitMask::op_Subtraction(BitMask,UInt32).0.arrayc8aa351a91a705be1462d4711470c40b589d09135c08d50b79a45acfa9e94d27\(to_integer(to_signed(0, 32))) := \BitMask::op_Subtraction(BitMask,UInt32).0.right\;
                        -- Initializing record fields to their defaults.
                        \BitMask::op_Subtraction(BitMask,UInt32).0.object77d16c4ef26cad24ef177b742166d622e968246a8b3c1e923c73e932760e2cc3\.\IsNull\ := false;
                        \BitMask::op_Subtraction(BitMask,UInt32).0.object77d16c4ef26cad24ef177b742166d622e968246a8b3c1e923c73e932760e2cc3\.\Size\ := to_unsigned(0, 16);
                        \BitMask::op_Subtraction(BitMask,UInt32).0.object77d16c4ef26cad24ef177b742166d622e968246a8b3c1e923c73e932760e2cc3\.\SegmentCount\ := to_unsigned(0, 16);
                        \BitMask::op_Subtraction(BitMask,UInt32).0.object77d16c4ef26cad24ef177b742166d622e968246a8b3c1e923c73e932760e2cc3\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\ <= \BitMask::op_Subtraction(BitMask,UInt32).0.object77d16c4ef26cad24ef177b742166d622e968246a8b3c1e923c73e932760e2cc3\;
                        \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\(0 to 0) <= \BitMask::op_Subtraction(BitMask,UInt32).0.arrayc8aa351a91a705be1462d4711470c40b589d09135c08d50b79a45acfa9e94d27\;
                        \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= \BitMask::op_Subtraction(BitMask,UInt32).0.left\.\Size\;
                        \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= true;
                        \BitMask::op_Subtraction(BitMask,UInt32).0._State\ := \BitMask::op_Subtraction(BitMask,UInt32).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Subtraction(BitMask,UInt32).0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        if (\BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\) then 
                            \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                            \BitMask::op_Subtraction(BitMask,UInt32).0.object77d16c4ef26cad24ef177b742166d622e968246a8b3c1e923c73e932760e2cc3\ := \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\;
                            \BitMask::op_Subtraction(BitMask,UInt32).0.arrayc8aa351a91a705be1462d4711470c40b589d09135c08d50b79a45acfa9e94d27\ := \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\(0 to 0);
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::op_Subtraction(BitMask,BitMask).left.parameter.Out.0\ <= \BitMask::op_Subtraction(BitMask,UInt32).0.left\;
                            \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::op_Subtraction(BitMask,BitMask).right.parameter.Out.0\ <= \BitMask::op_Subtraction(BitMask,UInt32).0.object77d16c4ef26cad24ef177b742166d622e968246a8b3c1e923c73e932760e2cc3\;
                            \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ <= true;
                            \BitMask::op_Subtraction(BitMask,UInt32).0._State\ := \BitMask::op_Subtraction(BitMask,UInt32).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Subtraction(BitMask,UInt32).0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ = \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::op_Subtraction(BitMask,BitMask)._Finished.0\) then 
                            \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ <= false;
                            \BitMask::op_Subtraction(BitMask,UInt32).0.return.0\ := \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::op_Subtraction(BitMask,BitMask).return.0\;
                            \BitMask::op_Subtraction(BitMask,UInt32).0.return\ <= \BitMask::op_Subtraction(BitMask,UInt32).0.return.0\;
                            \BitMask::op_Subtraction(BitMask,UInt32).0._State\ := \BitMask::op_Subtraction(BitMask,UInt32).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,System.UInt32).0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 state machine start
    \BitMask::op_Addition(BitMask,BitMask).0._StateMachine\: process (\Clock\) 
        Variable \BitMask::op_Addition(BitMask,BitMask).0._State\: \BitMask::op_Addition(BitMask,BitMask).0._States\ := \BitMask::op_Addition(BitMask,BitMask).0._State_0\;
        Variable \BitMask::op_Addition(BitMask,BitMask).0.left\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_Addition(BitMask,BitMask).0.right\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_Addition(BitMask,BitMask).0.flag\: boolean := false;
        Variable \BitMask::op_Addition(BitMask,BitMask).0.result\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_Addition(BitMask,BitMask).0.flag2\: boolean := false;
        Variable \BitMask::op_Addition(BitMask,BitMask).0.num\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.num2\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.array\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
        Variable \BitMask::op_Addition(BitMask,BitMask).0.num3\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.flag3\: boolean := false;
        Variable \BitMask::op_Addition(BitMask,BitMask).0.flag4\: boolean := false;
        Variable \BitMask::op_Addition(BitMask,BitMask).0.b\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.flag5\: boolean := false;
        Variable \BitMask::op_Addition(BitMask,BitMask).0.flag6\: boolean := false;
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.0\: boolean := false;
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.1\: boolean := false;
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.2\: boolean := false;
        Variable \BitMask::op_Addition(BitMask,BitMask).0.conditional634a6c6c4335747fbb3127d03ed2dabb2d062c45b344366ead52f18db6080904\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.3\: boolean := false;
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.4\: boolean := false;
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.5\: boolean := false;
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.6\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.7\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.8\: boolean := false;
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.9\: boolean := false;
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.10\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.11\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.12\: boolean := false;
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.13\: boolean := false;
        Variable \BitMask::op_Addition(BitMask,BitMask).0.conditionale434122820f41deb9aa7a0d1af32faf6cb55e904d124344b6c6dafef1d0a4000\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.conditionalab620eac6807dc6e4094d422af6311ede25245ae0b71988698e3f0d88867f131\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.conditional8b600d3c1f6fe3101e3ae23b08db358034ba82e520e35fd6640dd2e72d7ef7d5\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.14\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.15\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.16\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.17\: boolean := false;
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.18\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.19\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.20\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.21\: boolean := false;
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.22\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.23\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.24\: boolean := false;
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.25\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.26\: unsigned(15 downto 0) := to_unsigned(0, 16);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \BitMask::op_Addition(BitMask,BitMask).0._Finished\ <= false;
                \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 32));
                \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_0\;
                \BitMask::op_Addition(BitMask,BitMask).0.flag\ := false;
                \BitMask::op_Addition(BitMask,BitMask).0.flag2\ := false;
                \BitMask::op_Addition(BitMask,BitMask).0.num\ := to_unsigned(0, 16);
                \BitMask::op_Addition(BitMask,BitMask).0.num2\ := to_unsigned(0, 16);
                \BitMask::op_Addition(BitMask,BitMask).0.array\ := (others => to_unsigned(0, 32));
                \BitMask::op_Addition(BitMask,BitMask).0.num3\ := to_unsigned(0, 16);
                \BitMask::op_Addition(BitMask,BitMask).0.flag3\ := false;
                \BitMask::op_Addition(BitMask,BitMask).0.flag4\ := false;
                \BitMask::op_Addition(BitMask,BitMask).0.b\ := to_unsigned(0, 8);
                \BitMask::op_Addition(BitMask,BitMask).0.flag5\ := false;
                \BitMask::op_Addition(BitMask,BitMask).0.flag6\ := false;
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.0\ := false;
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.1\ := false;
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.2\ := false;
                \BitMask::op_Addition(BitMask,BitMask).0.conditional634a6c6c4335747fbb3127d03ed2dabb2d062c45b344366ead52f18db6080904\ := to_unsigned(0, 16);
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.3\ := false;
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.4\ := false;
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.5\ := false;
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.6\ := to_unsigned(0, 32);
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.7\ := to_unsigned(0, 32);
                \BitMask::op_Addition(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.8\ := false;
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.9\ := false;
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.10\ := to_unsigned(0, 32);
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.11\ := to_unsigned(0, 32);
                \BitMask::op_Addition(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.1\ := to_signed(0, 32);
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.12\ := false;
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.13\ := false;
                \BitMask::op_Addition(BitMask,BitMask).0.conditionale434122820f41deb9aa7a0d1af32faf6cb55e904d124344b6c6dafef1d0a4000\ := to_signed(0, 32);
                \BitMask::op_Addition(BitMask,BitMask).0.conditionalab620eac6807dc6e4094d422af6311ede25245ae0b71988698e3f0d88867f131\ := to_signed(0, 32);
                \BitMask::op_Addition(BitMask,BitMask).0.conditional8b600d3c1f6fe3101e3ae23b08db358034ba82e520e35fd6640dd2e72d7ef7d5\ := to_signed(0, 32);
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.14\ := to_signed(0, 32);
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.15\ := to_unsigned(0, 8);
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.16\ := to_unsigned(0, 8);
                \BitMask::op_Addition(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.2\ := to_signed(0, 32);
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.17\ := false;
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.18\ := to_unsigned(0, 32);
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.19\ := to_unsigned(0, 32);
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.20\ := to_signed(0, 32);
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.21\ := false;
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.22\ := to_unsigned(0, 16);
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.23\ := to_signed(0, 32);
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.24\ := false;
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.25\ := to_unsigned(0, 16);
                \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.26\ := to_unsigned(0, 16);
            else 
                case \BitMask::op_Addition(BitMask,BitMask).0._State\ is 
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\BitMask::op_Addition(BitMask,BitMask).0._Started\ = true) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\BitMask::op_Addition(BitMask,BitMask).0._Started\ = true) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._Finished\ <= true;
                        else 
                            \BitMask::op_Addition(BitMask,BitMask).0._Finished\ <= false;
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_2\ => 
                        \BitMask::op_Addition(BitMask,BitMask).0.left\ := \BitMask::op_Addition(BitMask,BitMask).0.left.parameter.In\;
                        \BitMask::op_Addition(BitMask,BitMask).0.right\ := \BitMask::op_Addition(BitMask,BitMask).0.right.parameter.In\;
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.0\ := \BitMask::op_Addition(BitMask,BitMask).0.left\.\SegmentCount\ = to_unsigned(0, 16);
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.1\ := \BitMask::op_Addition(BitMask,BitMask).0.right\.\SegmentCount\ = to_unsigned(0, 16);
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.2\ := \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.0\ or \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.1\;
                        \BitMask::op_Addition(BitMask,BitMask).0.flag\ := \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.2\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::op_Addition(BitMask,BitMask).0._State_4\ and ends in state \BitMask::op_Addition(BitMask,BitMask).0._State_4\.
                        --     * The false branch starts in state \BitMask::op_Addition(BitMask,BitMask).0._State_5\ and ends in state \BitMask::op_Addition(BitMask,BitMask).0._State_30\.
                        --     * Execution after either branch will continue in the following state: \BitMask::op_Addition(BitMask,BitMask).0._State_3\.

                        if (\BitMask::op_Addition(BitMask,BitMask).0.flag\) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_4\;
                        else 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_3\ => 
                        -- State after the if-else which was started in state \BitMask::op_Addition(BitMask,BitMask).0._State_2\.
                        \BitMask::op_Addition(BitMask,BitMask).0.return\ <= \BitMask::op_Addition(BitMask,BitMask).0.result\;
                        \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_4\ => 
                        -- True branch of the if-else started in state \BitMask::op_Addition(BitMask,BitMask).0._State_2\.
                        \BitMask::op_Addition(BitMask,BitMask).0.result\ := \BitMask::op_Addition(BitMask,BitMask).0.left\;
                        -- Going to the state after the if-else which was started in state \BitMask::op_Addition(BitMask,BitMask).0._State_2\.
                        if (\BitMask::op_Addition(BitMask,BitMask).0._State\ = \BitMask::op_Addition(BitMask,BitMask).0._State_4\) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_5\ => 
                        -- False branch of the if-else started in state \BitMask::op_Addition(BitMask,BitMask).0._State_2\.
                        \BitMask::op_Addition(BitMask,BitMask).0.flag2\ := False;
                        \BitMask::op_Addition(BitMask,BitMask).0.num\ := to_unsigned(0, 16);
                        \BitMask::op_Addition(BitMask,BitMask).0.num2\ := to_unsigned(0, 16);
                        \BitMask::op_Addition(BitMask,BitMask).0.array\ := (others => to_unsigned(0, 32));
                        \BitMask::op_Addition(BitMask,BitMask).0.num3\ := to_unsigned(0, 16);
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.3\ := \BitMask::op_Addition(BitMask,BitMask).0.left\.\Size\ > \BitMask::op_Addition(BitMask,BitMask).0.right\.\Size\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::op_Addition(BitMask,BitMask).0._State_7\ and ends in state \BitMask::op_Addition(BitMask,BitMask).0._State_7\.
                        --     * The false branch starts in state \BitMask::op_Addition(BitMask,BitMask).0._State_8\ and ends in state \BitMask::op_Addition(BitMask,BitMask).0._State_8\.
                        --     * Execution after either branch will continue in the following state: \BitMask::op_Addition(BitMask,BitMask).0._State_6\.

                        if (\BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.3\) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_7\;
                        else 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_6\ => 
                        -- State after the if-else which was started in state \BitMask::op_Addition(BitMask,BitMask).0._State_5\.
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.4\ := \BitMask::op_Addition(BitMask,BitMask).0.num3\ < \BitMask::op_Addition(BitMask,BitMask).0.conditional634a6c6c4335747fbb3127d03ed2dabb2d062c45b344366ead52f18db6080904\;
                        if (\BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.4\) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_9\;
                        else 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_10\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_7\ => 
                        -- True branch of the if-else started in state \BitMask::op_Addition(BitMask,BitMask).0._State_5\.
                        \BitMask::op_Addition(BitMask,BitMask).0.conditional634a6c6c4335747fbb3127d03ed2dabb2d062c45b344366ead52f18db6080904\ := \BitMask::op_Addition(BitMask,BitMask).0.left\.\Size\;
                        -- Going to the state after the if-else which was started in state \BitMask::op_Addition(BitMask,BitMask).0._State_5\.
                        if (\BitMask::op_Addition(BitMask,BitMask).0._State\ = \BitMask::op_Addition(BitMask,BitMask).0._State_7\) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_8\ => 
                        -- False branch of the if-else started in state \BitMask::op_Addition(BitMask,BitMask).0._State_5\.
                        \BitMask::op_Addition(BitMask,BitMask).0.conditional634a6c6c4335747fbb3127d03ed2dabb2d062c45b344366ead52f18db6080904\ := \BitMask::op_Addition(BitMask,BitMask).0.right\.\Size\;
                        -- Going to the state after the if-else which was started in state \BitMask::op_Addition(BitMask,BitMask).0._State_5\.
                        if (\BitMask::op_Addition(BitMask,BitMask).0._State\ = \BitMask::op_Addition(BitMask,BitMask).0._State_8\) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_9\ => 
                        -- Repeated state of the while loop which was started in state \BitMask::op_Addition(BitMask,BitMask).0._State_6\.
                        -- The while loop's condition:
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.5\ := \BitMask::op_Addition(BitMask,BitMask).0.num3\ < \BitMask::op_Addition(BitMask,BitMask).0.conditional634a6c6c4335747fbb3127d03ed2dabb2d062c45b344366ead52f18db6080904\;
                        if (\BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.5\) then 
                            \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.6\ := resize(shift_right(\BitMask::op_Addition(BitMask,BitMask).0.left\.\Segments\(to_integer(resize(signed(\BitMask::op_Addition(BitMask,BitMask).0.num\), 32))), to_integer(resize(signed(\BitMask::op_Addition(BitMask,BitMask).0.num2\), 32))), 32);
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_11\;
                        else 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_10\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_10\ => 
                        -- State after the while loop which was started in state \BitMask::op_Addition(BitMask,BitMask).0._State_6\.
                        -- Initializing record fields to their defaults.
                        \BitMask::op_Addition(BitMask,BitMask).0.result\.\IsNull\ := false;
                        \BitMask::op_Addition(BitMask,BitMask).0.result\.\Size\ := to_unsigned(0, 16);
                        \BitMask::op_Addition(BitMask,BitMask).0.result\.\SegmentCount\ := to_unsigned(0, 16);
                        \BitMask::op_Addition(BitMask,BitMask).0.result\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\ <= \BitMask::op_Addition(BitMask,BitMask).0.result\;
                        \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\ <= \BitMask::op_Addition(BitMask,BitMask).0.array\;
                        \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                        \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= true;
                        \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_30\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_11\ => 
                        -- Waiting for the result to appear in \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.7\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\BitMask::op_Addition(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_12\;
                            \BitMask::op_Addition(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \BitMask::op_Addition(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.0\ := \BitMask::op_Addition(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.7\ := \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.6\ mod to_unsigned(2, 32);
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_12\ => 
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.8\ := \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.7\ = to_unsigned(1, 32);
                        \BitMask::op_Addition(BitMask,BitMask).0.flag3\ := \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.8\;
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.9\ := \BitMask::op_Addition(BitMask,BitMask).0.num3\ < \BitMask::op_Addition(BitMask,BitMask).0.right\.\Size\;
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.10\ := resize(shift_right(\BitMask::op_Addition(BitMask,BitMask).0.right\.\Segments\(to_integer(resize(signed(\BitMask::op_Addition(BitMask,BitMask).0.num\), 32))), to_integer(resize(signed(\BitMask::op_Addition(BitMask,BitMask).0.num2\), 32))), 32);
                        \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_13\;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_13\ => 
                        -- Waiting for the result to appear in \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.11\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\BitMask::op_Addition(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.1\ >= to_signed(7, 32)) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_14\;
                            \BitMask::op_Addition(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.1\ := to_signed(0, 32);
                        else 
                            \BitMask::op_Addition(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.1\ := \BitMask::op_Addition(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.1\ + to_signed(1, 32);
                        end if;
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.11\ := \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.10\ mod to_unsigned(2, 32);
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_14\ => 
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.12\ := \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.11\ = to_unsigned(1, 32);
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.13\ := \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.9\ and \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.12\;
                        \BitMask::op_Addition(BitMask,BitMask).0.flag4\ := \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.13\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::op_Addition(BitMask,BitMask).0._State_16\ and ends in state \BitMask::op_Addition(BitMask,BitMask).0._State_16\.
                        --     * The false branch starts in state \BitMask::op_Addition(BitMask,BitMask).0._State_17\ and ends in state \BitMask::op_Addition(BitMask,BitMask).0._State_17\.
                        --     * Execution after either branch will continue in the following state: \BitMask::op_Addition(BitMask,BitMask).0._State_15\.

                        if (\BitMask::op_Addition(BitMask,BitMask).0.flag3\) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_16\;
                        else 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_17\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_15\ => 
                        -- State after the if-else which was started in state \BitMask::op_Addition(BitMask,BitMask).0._State_14\.

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::op_Addition(BitMask,BitMask).0._State_19\ and ends in state \BitMask::op_Addition(BitMask,BitMask).0._State_19\.
                        --     * The false branch starts in state \BitMask::op_Addition(BitMask,BitMask).0._State_20\ and ends in state \BitMask::op_Addition(BitMask,BitMask).0._State_20\.
                        --     * Execution after either branch will continue in the following state: \BitMask::op_Addition(BitMask,BitMask).0._State_18\.

                        if (\BitMask::op_Addition(BitMask,BitMask).0.flag4\) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_19\;
                        else 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_20\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_16\ => 
                        -- True branch of the if-else started in state \BitMask::op_Addition(BitMask,BitMask).0._State_14\.
                        \BitMask::op_Addition(BitMask,BitMask).0.conditionale434122820f41deb9aa7a0d1af32faf6cb55e904d124344b6c6dafef1d0a4000\ := to_signed(1, 32);
                        -- Going to the state after the if-else which was started in state \BitMask::op_Addition(BitMask,BitMask).0._State_14\.
                        if (\BitMask::op_Addition(BitMask,BitMask).0._State\ = \BitMask::op_Addition(BitMask,BitMask).0._State_16\) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_15\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_17\ => 
                        -- False branch of the if-else started in state \BitMask::op_Addition(BitMask,BitMask).0._State_14\.
                        \BitMask::op_Addition(BitMask,BitMask).0.conditionale434122820f41deb9aa7a0d1af32faf6cb55e904d124344b6c6dafef1d0a4000\ := to_signed(0, 32);
                        -- Going to the state after the if-else which was started in state \BitMask::op_Addition(BitMask,BitMask).0._State_14\.
                        if (\BitMask::op_Addition(BitMask,BitMask).0._State\ = \BitMask::op_Addition(BitMask,BitMask).0._State_17\) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_15\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_18\ => 
                        -- State after the if-else which was started in state \BitMask::op_Addition(BitMask,BitMask).0._State_15\.

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::op_Addition(BitMask,BitMask).0._State_22\ and ends in state \BitMask::op_Addition(BitMask,BitMask).0._State_22\.
                        --     * The false branch starts in state \BitMask::op_Addition(BitMask,BitMask).0._State_23\ and ends in state \BitMask::op_Addition(BitMask,BitMask).0._State_23\.
                        --     * Execution after either branch will continue in the following state: \BitMask::op_Addition(BitMask,BitMask).0._State_21\.

                        if (\BitMask::op_Addition(BitMask,BitMask).0.flag2\) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_22\;
                        else 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_23\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_19\ => 
                        -- True branch of the if-else started in state \BitMask::op_Addition(BitMask,BitMask).0._State_15\.
                        \BitMask::op_Addition(BitMask,BitMask).0.conditionalab620eac6807dc6e4094d422af6311ede25245ae0b71988698e3f0d88867f131\ := to_signed(1, 32);
                        -- Going to the state after the if-else which was started in state \BitMask::op_Addition(BitMask,BitMask).0._State_15\.
                        if (\BitMask::op_Addition(BitMask,BitMask).0._State\ = \BitMask::op_Addition(BitMask,BitMask).0._State_19\) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_18\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_20\ => 
                        -- False branch of the if-else started in state \BitMask::op_Addition(BitMask,BitMask).0._State_15\.
                        \BitMask::op_Addition(BitMask,BitMask).0.conditionalab620eac6807dc6e4094d422af6311ede25245ae0b71988698e3f0d88867f131\ := to_signed(0, 32);
                        -- Going to the state after the if-else which was started in state \BitMask::op_Addition(BitMask,BitMask).0._State_15\.
                        if (\BitMask::op_Addition(BitMask,BitMask).0._State\ = \BitMask::op_Addition(BitMask,BitMask).0._State_20\) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_18\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_21\ => 
                        -- State after the if-else which was started in state \BitMask::op_Addition(BitMask,BitMask).0._State_18\.
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.14\ := \BitMask::op_Addition(BitMask,BitMask).0.conditionale434122820f41deb9aa7a0d1af32faf6cb55e904d124344b6c6dafef1d0a4000\ + \BitMask::op_Addition(BitMask,BitMask).0.conditionalab620eac6807dc6e4094d422af6311ede25245ae0b71988698e3f0d88867f131\;
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.15\ := resize(unsigned(\BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.14\ + \BitMask::op_Addition(BitMask,BitMask).0.conditional8b600d3c1f6fe3101e3ae23b08db358034ba82e520e35fd6640dd2e72d7ef7d5\), 8);
                        \BitMask::op_Addition(BitMask,BitMask).0.b\ := (\BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.15\);
                        \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_24\;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_22\ => 
                        -- True branch of the if-else started in state \BitMask::op_Addition(BitMask,BitMask).0._State_18\.
                        \BitMask::op_Addition(BitMask,BitMask).0.conditional8b600d3c1f6fe3101e3ae23b08db358034ba82e520e35fd6640dd2e72d7ef7d5\ := to_signed(1, 32);
                        -- Going to the state after the if-else which was started in state \BitMask::op_Addition(BitMask,BitMask).0._State_18\.
                        if (\BitMask::op_Addition(BitMask,BitMask).0._State\ = \BitMask::op_Addition(BitMask,BitMask).0._State_22\) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_21\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_23\ => 
                        -- False branch of the if-else started in state \BitMask::op_Addition(BitMask,BitMask).0._State_18\.
                        \BitMask::op_Addition(BitMask,BitMask).0.conditional8b600d3c1f6fe3101e3ae23b08db358034ba82e520e35fd6640dd2e72d7ef7d5\ := to_signed(0, 32);
                        -- Going to the state after the if-else which was started in state \BitMask::op_Addition(BitMask,BitMask).0._State_18\.
                        if (\BitMask::op_Addition(BitMask,BitMask).0._State\ = \BitMask::op_Addition(BitMask,BitMask).0._State_23\) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_21\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_24\ => 
                        -- Waiting for the result to appear in \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.16\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\BitMask::op_Addition(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.2\ >= to_signed(7, 32)) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_25\;
                            \BitMask::op_Addition(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.2\ := to_signed(0, 32);
                        else 
                            \BitMask::op_Addition(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.2\ := \BitMask::op_Addition(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.2\ + to_signed(1, 32);
                        end if;
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.16\ := \BitMask::op_Addition(BitMask,BitMask).0.b\ mod to_unsigned(2, 8);
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_25\ => 
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.17\ := \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.16\ = to_unsigned(1, 8);
                        \BitMask::op_Addition(BitMask,BitMask).0.flag5\ := \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.17\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::op_Addition(BitMask,BitMask).0._State_27\ and ends in state \BitMask::op_Addition(BitMask,BitMask).0._State_27\.
                        --     * Execution after either branch will continue in the following state: \BitMask::op_Addition(BitMask,BitMask).0._State_26\.

                        if (\BitMask::op_Addition(BitMask,BitMask).0.flag5\) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_27\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_26\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_26\ => 
                        -- State after the if-else which was started in state \BitMask::op_Addition(BitMask,BitMask).0._State_25\.
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.20\ := resize(signed(shift_right(\BitMask::op_Addition(BitMask,BitMask).0.b\, to_integer(to_signed(1, 32)))), 32);
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.21\ := \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.20\ = to_signed(1, 32);
                        \BitMask::op_Addition(BitMask,BitMask).0.flag2\ := \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.21\;
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.22\ := \BitMask::op_Addition(BitMask,BitMask).0.num2\ + to_unsigned(1, 16);
                        \BitMask::op_Addition(BitMask,BitMask).0.num2\ := \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.22\;
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.23\ := resize(signed(shift_right(\BitMask::op_Addition(BitMask,BitMask).0.num2\, to_integer(to_signed(5, 32)))), 32);
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.24\ := \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.23\ = to_signed(1, 32);
                        \BitMask::op_Addition(BitMask,BitMask).0.flag6\ := \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.24\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::op_Addition(BitMask,BitMask).0._State_29\ and ends in state \BitMask::op_Addition(BitMask,BitMask).0._State_29\.
                        --     * Execution after either branch will continue in the following state: \BitMask::op_Addition(BitMask,BitMask).0._State_28\.

                        if (\BitMask::op_Addition(BitMask,BitMask).0.flag6\) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_29\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_28\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.5
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_27\ => 
                        -- True branch of the if-else started in state \BitMask::op_Addition(BitMask,BitMask).0._State_25\.
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.18\ := resize(shift_left(to_unsigned(1, 32), to_integer(resize(signed(\BitMask::op_Addition(BitMask,BitMask).0.num2\), 32))), 32);
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.19\ := \BitMask::op_Addition(BitMask,BitMask).0.array\(to_integer(resize(signed(\BitMask::op_Addition(BitMask,BitMask).0.num\), 32))) + \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.18\;
                        \BitMask::op_Addition(BitMask,BitMask).0.array\(to_integer(resize(signed(\BitMask::op_Addition(BitMask,BitMask).0.num\), 32))) := \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.19\;
                        -- Going to the state after the if-else which was started in state \BitMask::op_Addition(BitMask,BitMask).0._State_25\.
                        if (\BitMask::op_Addition(BitMask,BitMask).0._State\ = \BitMask::op_Addition(BitMask,BitMask).0._State_27\) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_26\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_28\ => 
                        -- State after the if-else which was started in state \BitMask::op_Addition(BitMask,BitMask).0._State_26\.
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.26\ := \BitMask::op_Addition(BitMask,BitMask).0.num3\ + to_unsigned(1, 16);
                        \BitMask::op_Addition(BitMask,BitMask).0.num3\ := \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.26\;
                        -- Returning to the repeated state of the while loop which was started in state \BitMask::op_Addition(BitMask,BitMask).0._State_6\ if the loop wasn't exited with a state change.
                        if (\BitMask::op_Addition(BitMask,BitMask).0._State\ = \BitMask::op_Addition(BitMask,BitMask).0._State_28\) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_9\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_29\ => 
                        -- True branch of the if-else started in state \BitMask::op_Addition(BitMask,BitMask).0._State_26\.
                        \BitMask::op_Addition(BitMask,BitMask).0.num2\ := to_unsigned(0, 16);
                        \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.25\ := \BitMask::op_Addition(BitMask,BitMask).0.num\ + to_unsigned(1, 16);
                        \BitMask::op_Addition(BitMask,BitMask).0.num\ := \BitMask::op_Addition(BitMask,BitMask).0.binaryOperationResult.25\;
                        -- Going to the state after the if-else which was started in state \BitMask::op_Addition(BitMask,BitMask).0._State_26\.
                        if (\BitMask::op_Addition(BitMask,BitMask).0._State\ = \BitMask::op_Addition(BitMask,BitMask).0._State_29\) then 
                            \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_28\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_Addition(BitMask,BitMask).0._State_30\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        if (\BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\) then 
                            \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                            \BitMask::op_Addition(BitMask,BitMask).0.result\ := \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\;
                            \BitMask::op_Addition(BitMask,BitMask).0.array\ := \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\;
                            -- Going to the state after the if-else which was started in state \BitMask::op_Addition(BitMask,BitMask).0._State_2\.
                            if (\BitMask::op_Addition(BitMask,BitMask).0._State\ = \BitMask::op_Addition(BitMask,BitMask).0._State_30\) then 
                                \BitMask::op_Addition(BitMask,BitMask).0._State\ := \BitMask::op_Addition(BitMask,BitMask).0._State_3\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 state machine start
    \BitMask::op_Subtraction(BitMask,BitMask).0._StateMachine\: process (\Clock\) 
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0._State\: \BitMask::op_Subtraction(BitMask,BitMask).0._States\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_0\;
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.left\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.right\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.flag\: boolean := false;
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.result\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.flag2\: boolean := false;
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.num\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.num2\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.array\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.num3\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.flag3\: boolean := false;
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.flag4\: boolean := false;
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.b\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.flag5\: boolean := false;
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.flag6\: boolean := false;
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.0\: boolean := false;
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.1\: boolean := false;
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.2\: boolean := false;
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.conditional634a6c6c4335747fbb3127d03ed2dabb2d062c45b344366ead52f18db6080904\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.3\: boolean := false;
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.4\: boolean := false;
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.5\: boolean := false;
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.6\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.7\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.8\: boolean := false;
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.9\: boolean := false;
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.10\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.11\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.12\: boolean := false;
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.13\: boolean := false;
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.conditionale434122820f41deb9aa7a0d1af32faf6cb55e904d124344b6c6dafef1d0a4000\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.conditionalab620eac6807dc6e4094d422af6311ede25245ae0b71988698e3f0d88867f131\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.conditional8b600d3c1f6fe3101e3ae23b08db358034ba82e520e35fd6640dd2e72d7ef7d5\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.14\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.15\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.16\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.17\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.18\: boolean := false;
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.19\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.20\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.21\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.22\: boolean := false;
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.23\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.24\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.25\: boolean := false;
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.26\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.27\: unsigned(15 downto 0) := to_unsigned(0, 16);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \BitMask::op_Subtraction(BitMask,BitMask).0._Finished\ <= false;
                \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 32));
                \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_0\;
                \BitMask::op_Subtraction(BitMask,BitMask).0.flag\ := false;
                \BitMask::op_Subtraction(BitMask,BitMask).0.flag2\ := false;
                \BitMask::op_Subtraction(BitMask,BitMask).0.num\ := to_unsigned(0, 16);
                \BitMask::op_Subtraction(BitMask,BitMask).0.num2\ := to_unsigned(0, 16);
                \BitMask::op_Subtraction(BitMask,BitMask).0.array\ := (others => to_unsigned(0, 32));
                \BitMask::op_Subtraction(BitMask,BitMask).0.num3\ := to_unsigned(0, 16);
                \BitMask::op_Subtraction(BitMask,BitMask).0.flag3\ := false;
                \BitMask::op_Subtraction(BitMask,BitMask).0.flag4\ := false;
                \BitMask::op_Subtraction(BitMask,BitMask).0.b\ := to_unsigned(0, 8);
                \BitMask::op_Subtraction(BitMask,BitMask).0.flag5\ := false;
                \BitMask::op_Subtraction(BitMask,BitMask).0.flag6\ := false;
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.0\ := false;
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.1\ := false;
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.2\ := false;
                \BitMask::op_Subtraction(BitMask,BitMask).0.conditional634a6c6c4335747fbb3127d03ed2dabb2d062c45b344366ead52f18db6080904\ := to_unsigned(0, 16);
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.3\ := false;
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.4\ := false;
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.5\ := false;
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.6\ := to_unsigned(0, 32);
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.7\ := to_unsigned(0, 32);
                \BitMask::op_Subtraction(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.8\ := false;
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.9\ := false;
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.10\ := to_unsigned(0, 32);
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.11\ := to_unsigned(0, 32);
                \BitMask::op_Subtraction(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.1\ := to_signed(0, 32);
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.12\ := false;
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.13\ := false;
                \BitMask::op_Subtraction(BitMask,BitMask).0.conditionale434122820f41deb9aa7a0d1af32faf6cb55e904d124344b6c6dafef1d0a4000\ := to_signed(0, 32);
                \BitMask::op_Subtraction(BitMask,BitMask).0.conditionalab620eac6807dc6e4094d422af6311ede25245ae0b71988698e3f0d88867f131\ := to_signed(0, 32);
                \BitMask::op_Subtraction(BitMask,BitMask).0.conditional8b600d3c1f6fe3101e3ae23b08db358034ba82e520e35fd6640dd2e72d7ef7d5\ := to_signed(0, 32);
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.14\ := to_signed(0, 32);
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.15\ := to_signed(0, 32);
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.16\ := to_unsigned(0, 8);
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.17\ := to_unsigned(0, 8);
                \BitMask::op_Subtraction(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.2\ := to_signed(0, 32);
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.18\ := false;
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.19\ := to_unsigned(0, 32);
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.20\ := to_unsigned(0, 32);
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.21\ := to_signed(0, 32);
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.22\ := false;
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.23\ := to_unsigned(0, 16);
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.24\ := to_signed(0, 32);
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.25\ := false;
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.26\ := to_unsigned(0, 16);
                \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.27\ := to_unsigned(0, 16);
            else 
                case \BitMask::op_Subtraction(BitMask,BitMask).0._State\ is 
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\BitMask::op_Subtraction(BitMask,BitMask).0._Started\ = true) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\BitMask::op_Subtraction(BitMask,BitMask).0._Started\ = true) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._Finished\ <= true;
                        else 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._Finished\ <= false;
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_2\ => 
                        \BitMask::op_Subtraction(BitMask,BitMask).0.left\ := \BitMask::op_Subtraction(BitMask,BitMask).0.left.parameter.In\;
                        \BitMask::op_Subtraction(BitMask,BitMask).0.right\ := \BitMask::op_Subtraction(BitMask,BitMask).0.right.parameter.In\;
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.0\ := \BitMask::op_Subtraction(BitMask,BitMask).0.left\.\SegmentCount\ = to_unsigned(0, 16);
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.1\ := \BitMask::op_Subtraction(BitMask,BitMask).0.right\.\SegmentCount\ = to_unsigned(0, 16);
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.2\ := \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.0\ or \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.1\;
                        \BitMask::op_Subtraction(BitMask,BitMask).0.flag\ := \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.2\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_4\ and ends in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_4\.
                        --     * The false branch starts in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_5\ and ends in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_30\.
                        --     * Execution after either branch will continue in the following state: \BitMask::op_Subtraction(BitMask,BitMask).0._State_3\.

                        if (\BitMask::op_Subtraction(BitMask,BitMask).0.flag\) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_4\;
                        else 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_3\ => 
                        -- State after the if-else which was started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_2\.
                        \BitMask::op_Subtraction(BitMask,BitMask).0.return\ <= \BitMask::op_Subtraction(BitMask,BitMask).0.result\;
                        \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_4\ => 
                        -- True branch of the if-else started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_2\.
                        \BitMask::op_Subtraction(BitMask,BitMask).0.result\ := \BitMask::op_Subtraction(BitMask,BitMask).0.left\;
                        -- Going to the state after the if-else which was started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_2\.
                        if (\BitMask::op_Subtraction(BitMask,BitMask).0._State\ = \BitMask::op_Subtraction(BitMask,BitMask).0._State_4\) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_5\ => 
                        -- False branch of the if-else started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_2\.
                        \BitMask::op_Subtraction(BitMask,BitMask).0.flag2\ := False;
                        \BitMask::op_Subtraction(BitMask,BitMask).0.num\ := to_unsigned(0, 16);
                        \BitMask::op_Subtraction(BitMask,BitMask).0.num2\ := to_unsigned(0, 16);
                        \BitMask::op_Subtraction(BitMask,BitMask).0.array\ := (others => to_unsigned(0, 32));
                        \BitMask::op_Subtraction(BitMask,BitMask).0.num3\ := to_unsigned(0, 16);
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.3\ := \BitMask::op_Subtraction(BitMask,BitMask).0.left\.\Size\ > \BitMask::op_Subtraction(BitMask,BitMask).0.right\.\Size\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_7\ and ends in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_7\.
                        --     * The false branch starts in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_8\ and ends in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_8\.
                        --     * Execution after either branch will continue in the following state: \BitMask::op_Subtraction(BitMask,BitMask).0._State_6\.

                        if (\BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.3\) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_7\;
                        else 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_6\ => 
                        -- State after the if-else which was started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_5\.
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.4\ := \BitMask::op_Subtraction(BitMask,BitMask).0.num3\ < \BitMask::op_Subtraction(BitMask,BitMask).0.conditional634a6c6c4335747fbb3127d03ed2dabb2d062c45b344366ead52f18db6080904\;
                        if (\BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.4\) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_9\;
                        else 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_10\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_7\ => 
                        -- True branch of the if-else started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_5\.
                        \BitMask::op_Subtraction(BitMask,BitMask).0.conditional634a6c6c4335747fbb3127d03ed2dabb2d062c45b344366ead52f18db6080904\ := \BitMask::op_Subtraction(BitMask,BitMask).0.left\.\Size\;
                        -- Going to the state after the if-else which was started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_5\.
                        if (\BitMask::op_Subtraction(BitMask,BitMask).0._State\ = \BitMask::op_Subtraction(BitMask,BitMask).0._State_7\) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_8\ => 
                        -- False branch of the if-else started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_5\.
                        \BitMask::op_Subtraction(BitMask,BitMask).0.conditional634a6c6c4335747fbb3127d03ed2dabb2d062c45b344366ead52f18db6080904\ := \BitMask::op_Subtraction(BitMask,BitMask).0.right\.\Size\;
                        -- Going to the state after the if-else which was started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_5\.
                        if (\BitMask::op_Subtraction(BitMask,BitMask).0._State\ = \BitMask::op_Subtraction(BitMask,BitMask).0._State_8\) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_9\ => 
                        -- Repeated state of the while loop which was started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_6\.
                        -- The while loop's condition:
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.5\ := \BitMask::op_Subtraction(BitMask,BitMask).0.num3\ < \BitMask::op_Subtraction(BitMask,BitMask).0.conditional634a6c6c4335747fbb3127d03ed2dabb2d062c45b344366ead52f18db6080904\;
                        if (\BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.5\) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.6\ := resize(shift_right(\BitMask::op_Subtraction(BitMask,BitMask).0.left\.\Segments\(to_integer(resize(signed(\BitMask::op_Subtraction(BitMask,BitMask).0.num\), 32))), to_integer(resize(signed(\BitMask::op_Subtraction(BitMask,BitMask).0.num2\), 32))), 32);
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_11\;
                        else 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_10\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_10\ => 
                        -- State after the while loop which was started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_6\.
                        -- Initializing record fields to their defaults.
                        \BitMask::op_Subtraction(BitMask,BitMask).0.result\.\IsNull\ := false;
                        \BitMask::op_Subtraction(BitMask,BitMask).0.result\.\Size\ := to_unsigned(0, 16);
                        \BitMask::op_Subtraction(BitMask,BitMask).0.result\.\SegmentCount\ := to_unsigned(0, 16);
                        \BitMask::op_Subtraction(BitMask,BitMask).0.result\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\ <= \BitMask::op_Subtraction(BitMask,BitMask).0.result\;
                        \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\ <= \BitMask::op_Subtraction(BitMask,BitMask).0.array\;
                        \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                        \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= true;
                        \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_30\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_11\ => 
                        -- Waiting for the result to appear in \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.7\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\BitMask::op_Subtraction(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_12\;
                            \BitMask::op_Subtraction(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \BitMask::op_Subtraction(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.0\ := \BitMask::op_Subtraction(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.7\ := \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.6\ mod to_unsigned(2, 32);
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_12\ => 
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.8\ := \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.7\ = to_unsigned(1, 32);
                        \BitMask::op_Subtraction(BitMask,BitMask).0.flag3\ := \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.8\;
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.9\ := \BitMask::op_Subtraction(BitMask,BitMask).0.num3\ < \BitMask::op_Subtraction(BitMask,BitMask).0.right\.\Size\;
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.10\ := resize(shift_right(\BitMask::op_Subtraction(BitMask,BitMask).0.right\.\Segments\(to_integer(resize(signed(\BitMask::op_Subtraction(BitMask,BitMask).0.num\), 32))), to_integer(resize(signed(\BitMask::op_Subtraction(BitMask,BitMask).0.num2\), 32))), 32);
                        \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_13\;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_13\ => 
                        -- Waiting for the result to appear in \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.11\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\BitMask::op_Subtraction(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.1\ >= to_signed(7, 32)) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_14\;
                            \BitMask::op_Subtraction(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.1\ := to_signed(0, 32);
                        else 
                            \BitMask::op_Subtraction(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.1\ := \BitMask::op_Subtraction(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.1\ + to_signed(1, 32);
                        end if;
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.11\ := \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.10\ mod to_unsigned(2, 32);
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_14\ => 
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.12\ := \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.11\ = to_unsigned(1, 32);
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.13\ := \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.9\ and \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.12\;
                        \BitMask::op_Subtraction(BitMask,BitMask).0.flag4\ := \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.13\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_16\ and ends in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_16\.
                        --     * The false branch starts in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_17\ and ends in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_17\.
                        --     * Execution after either branch will continue in the following state: \BitMask::op_Subtraction(BitMask,BitMask).0._State_15\.

                        if (\BitMask::op_Subtraction(BitMask,BitMask).0.flag3\) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_16\;
                        else 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_17\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_15\ => 
                        -- State after the if-else which was started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_14\.

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_19\ and ends in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_19\.
                        --     * The false branch starts in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_20\ and ends in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_20\.
                        --     * Execution after either branch will continue in the following state: \BitMask::op_Subtraction(BitMask,BitMask).0._State_18\.

                        if (\BitMask::op_Subtraction(BitMask,BitMask).0.flag4\) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_19\;
                        else 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_20\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_16\ => 
                        -- True branch of the if-else started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_14\.
                        \BitMask::op_Subtraction(BitMask,BitMask).0.conditionale434122820f41deb9aa7a0d1af32faf6cb55e904d124344b6c6dafef1d0a4000\ := to_signed(1, 32);
                        -- Going to the state after the if-else which was started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_14\.
                        if (\BitMask::op_Subtraction(BitMask,BitMask).0._State\ = \BitMask::op_Subtraction(BitMask,BitMask).0._State_16\) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_15\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_17\ => 
                        -- False branch of the if-else started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_14\.
                        \BitMask::op_Subtraction(BitMask,BitMask).0.conditionale434122820f41deb9aa7a0d1af32faf6cb55e904d124344b6c6dafef1d0a4000\ := to_signed(0, 32);
                        -- Going to the state after the if-else which was started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_14\.
                        if (\BitMask::op_Subtraction(BitMask,BitMask).0._State\ = \BitMask::op_Subtraction(BitMask,BitMask).0._State_17\) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_15\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_18\ => 
                        -- State after the if-else which was started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_15\.

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_22\ and ends in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_22\.
                        --     * The false branch starts in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_23\ and ends in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_23\.
                        --     * Execution after either branch will continue in the following state: \BitMask::op_Subtraction(BitMask,BitMask).0._State_21\.

                        if (\BitMask::op_Subtraction(BitMask,BitMask).0.flag2\) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_22\;
                        else 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_23\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_19\ => 
                        -- True branch of the if-else started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_15\.
                        \BitMask::op_Subtraction(BitMask,BitMask).0.conditionalab620eac6807dc6e4094d422af6311ede25245ae0b71988698e3f0d88867f131\ := to_signed(1, 32);
                        -- Going to the state after the if-else which was started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_15\.
                        if (\BitMask::op_Subtraction(BitMask,BitMask).0._State\ = \BitMask::op_Subtraction(BitMask,BitMask).0._State_19\) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_18\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_20\ => 
                        -- False branch of the if-else started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_15\.
                        \BitMask::op_Subtraction(BitMask,BitMask).0.conditionalab620eac6807dc6e4094d422af6311ede25245ae0b71988698e3f0d88867f131\ := to_signed(0, 32);
                        -- Going to the state after the if-else which was started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_15\.
                        if (\BitMask::op_Subtraction(BitMask,BitMask).0._State\ = \BitMask::op_Subtraction(BitMask,BitMask).0._State_20\) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_18\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_21\ => 
                        -- State after the if-else which was started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_18\.
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.14\ := to_signed(2, 32) + \BitMask::op_Subtraction(BitMask,BitMask).0.conditionale434122820f41deb9aa7a0d1af32faf6cb55e904d124344b6c6dafef1d0a4000\;
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.15\ := \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.14\ - \BitMask::op_Subtraction(BitMask,BitMask).0.conditionalab620eac6807dc6e4094d422af6311ede25245ae0b71988698e3f0d88867f131\;
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.16\ := resize(unsigned(\BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.15\ - \BitMask::op_Subtraction(BitMask,BitMask).0.conditional8b600d3c1f6fe3101e3ae23b08db358034ba82e520e35fd6640dd2e72d7ef7d5\), 8);
                        \BitMask::op_Subtraction(BitMask,BitMask).0.b\ := (\BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.16\);
                        \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_24\;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_22\ => 
                        -- True branch of the if-else started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_18\.
                        \BitMask::op_Subtraction(BitMask,BitMask).0.conditional8b600d3c1f6fe3101e3ae23b08db358034ba82e520e35fd6640dd2e72d7ef7d5\ := to_signed(1, 32);
                        -- Going to the state after the if-else which was started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_18\.
                        if (\BitMask::op_Subtraction(BitMask,BitMask).0._State\ = \BitMask::op_Subtraction(BitMask,BitMask).0._State_22\) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_21\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_23\ => 
                        -- False branch of the if-else started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_18\.
                        \BitMask::op_Subtraction(BitMask,BitMask).0.conditional8b600d3c1f6fe3101e3ae23b08db358034ba82e520e35fd6640dd2e72d7ef7d5\ := to_signed(0, 32);
                        -- Going to the state after the if-else which was started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_18\.
                        if (\BitMask::op_Subtraction(BitMask,BitMask).0._State\ = \BitMask::op_Subtraction(BitMask,BitMask).0._State_23\) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_21\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_24\ => 
                        -- Waiting for the result to appear in \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.17\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\BitMask::op_Subtraction(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.2\ >= to_signed(7, 32)) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_25\;
                            \BitMask::op_Subtraction(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.2\ := to_signed(0, 32);
                        else 
                            \BitMask::op_Subtraction(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.2\ := \BitMask::op_Subtraction(BitMask,BitMask).0.clockCyclesWaitedForBinaryOperationResult.2\ + to_signed(1, 32);
                        end if;
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.17\ := \BitMask::op_Subtraction(BitMask,BitMask).0.b\ mod to_unsigned(2, 8);
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_25\ => 
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.18\ := \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.17\ = to_unsigned(1, 8);
                        \BitMask::op_Subtraction(BitMask,BitMask).0.flag5\ := \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.18\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_27\ and ends in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_27\.
                        --     * Execution after either branch will continue in the following state: \BitMask::op_Subtraction(BitMask,BitMask).0._State_26\.

                        if (\BitMask::op_Subtraction(BitMask,BitMask).0.flag5\) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_27\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_26\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_26\ => 
                        -- State after the if-else which was started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_25\.
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.21\ := resize(signed(shift_right(\BitMask::op_Subtraction(BitMask,BitMask).0.b\, to_integer(to_signed(1, 32)))), 32);
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.22\ := \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.21\ = to_signed(0, 32);
                        \BitMask::op_Subtraction(BitMask,BitMask).0.flag2\ := \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.22\;
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.23\ := \BitMask::op_Subtraction(BitMask,BitMask).0.num2\ + to_unsigned(1, 16);
                        \BitMask::op_Subtraction(BitMask,BitMask).0.num2\ := \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.23\;
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.24\ := resize(signed(shift_right(\BitMask::op_Subtraction(BitMask,BitMask).0.num2\, to_integer(to_signed(5, 32)))), 32);
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.25\ := \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.24\ = to_signed(1, 32);
                        \BitMask::op_Subtraction(BitMask,BitMask).0.flag6\ := \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.25\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_29\ and ends in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_29\.
                        --     * Execution after either branch will continue in the following state: \BitMask::op_Subtraction(BitMask,BitMask).0._State_28\.

                        if (\BitMask::op_Subtraction(BitMask,BitMask).0.flag6\) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_29\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_28\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.5
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_27\ => 
                        -- True branch of the if-else started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_25\.
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.19\ := resize(shift_left(to_unsigned(1, 32), to_integer(resize(signed(\BitMask::op_Subtraction(BitMask,BitMask).0.num2\), 32))), 32);
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.20\ := \BitMask::op_Subtraction(BitMask,BitMask).0.array\(to_integer(resize(signed(\BitMask::op_Subtraction(BitMask,BitMask).0.num\), 32))) + \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.19\;
                        \BitMask::op_Subtraction(BitMask,BitMask).0.array\(to_integer(resize(signed(\BitMask::op_Subtraction(BitMask,BitMask).0.num\), 32))) := \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.20\;
                        -- Going to the state after the if-else which was started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_25\.
                        if (\BitMask::op_Subtraction(BitMask,BitMask).0._State\ = \BitMask::op_Subtraction(BitMask,BitMask).0._State_27\) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_26\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_28\ => 
                        -- State after the if-else which was started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_26\.
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.27\ := \BitMask::op_Subtraction(BitMask,BitMask).0.num3\ + to_unsigned(1, 16);
                        \BitMask::op_Subtraction(BitMask,BitMask).0.num3\ := \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.27\;
                        -- Returning to the repeated state of the while loop which was started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_6\ if the loop wasn't exited with a state change.
                        if (\BitMask::op_Subtraction(BitMask,BitMask).0._State\ = \BitMask::op_Subtraction(BitMask,BitMask).0._State_28\) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_9\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_29\ => 
                        -- True branch of the if-else started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_26\.
                        \BitMask::op_Subtraction(BitMask,BitMask).0.num2\ := to_unsigned(0, 16);
                        \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.26\ := \BitMask::op_Subtraction(BitMask,BitMask).0.num\ + to_unsigned(1, 16);
                        \BitMask::op_Subtraction(BitMask,BitMask).0.num\ := \BitMask::op_Subtraction(BitMask,BitMask).0.binaryOperationResult.26\;
                        -- Going to the state after the if-else which was started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_26\.
                        if (\BitMask::op_Subtraction(BitMask,BitMask).0._State\ = \BitMask::op_Subtraction(BitMask,BitMask).0._State_29\) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_28\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_Subtraction(BitMask,BitMask).0._State_30\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        if (\BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                            \BitMask::op_Subtraction(BitMask,BitMask).0.result\ := \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\;
                            \BitMask::op_Subtraction(BitMask,BitMask).0.array\ := \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\;
                            -- Going to the state after the if-else which was started in state \BitMask::op_Subtraction(BitMask,BitMask).0._State_2\.
                            if (\BitMask::op_Subtraction(BitMask,BitMask).0._State\ = \BitMask::op_Subtraction(BitMask,BitMask).0._State_30\) then 
                                \BitMask::op_Subtraction(BitMask,BitMask).0._State\ := \BitMask::op_Subtraction(BitMask,BitMask).0._State_3\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseOr(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 state machine start
    \BitMask::op_BitwiseOr(BitMask,BitMask).0._StateMachine\: process (\Clock\) 
        Variable \BitMask::op_BitwiseOr(BitMask,BitMask).0._State\: \BitMask::op_BitwiseOr(BitMask,BitMask).0._States\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_0\;
        Variable \BitMask::op_BitwiseOr(BitMask,BitMask).0.left\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_BitwiseOr(BitMask,BitMask).0.right\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_BitwiseOr(BitMask,BitMask).0.flag\: boolean := false;
        Variable \BitMask::op_BitwiseOr(BitMask,BitMask).0.result\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_BitwiseOr(BitMask,BitMask).0.array\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
        Variable \BitMask::op_BitwiseOr(BitMask,BitMask).0.num\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_BitwiseOr(BitMask,BitMask).0.binaryOperationResult.0\: boolean := false;
        Variable \BitMask::op_BitwiseOr(BitMask,BitMask).0.binaryOperationResult.1\: boolean := false;
        Variable \BitMask::op_BitwiseOr(BitMask,BitMask).0.binaryOperationResult.2\: boolean := false;
        Variable \BitMask::op_BitwiseOr(BitMask,BitMask).0.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_BitwiseOr(BitMask,BitMask).0.binaryOperationResult.4\: unsigned(15 downto 0) := to_unsigned(0, 16);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \BitMask::op_BitwiseOr(BitMask,BitMask).0._Finished\ <= false;
                \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\ <= false;
                \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= false;
                \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 32));
                \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                \BitMask::op_BitwiseOr(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_0\;
                \BitMask::op_BitwiseOr(BitMask,BitMask).0.flag\ := false;
                \BitMask::op_BitwiseOr(BitMask,BitMask).0.array\ := (others => to_unsigned(0, 32));
                \BitMask::op_BitwiseOr(BitMask,BitMask).0.num\ := to_unsigned(0, 16);
                \BitMask::op_BitwiseOr(BitMask,BitMask).0.binaryOperationResult.0\ := false;
                \BitMask::op_BitwiseOr(BitMask,BitMask).0.binaryOperationResult.1\ := false;
                \BitMask::op_BitwiseOr(BitMask,BitMask).0.binaryOperationResult.2\ := false;
                \BitMask::op_BitwiseOr(BitMask,BitMask).0.binaryOperationResult.3\ := to_unsigned(0, 32);
                \BitMask::op_BitwiseOr(BitMask,BitMask).0.binaryOperationResult.4\ := to_unsigned(0, 16);
            else 
                case \BitMask::op_BitwiseOr(BitMask,BitMask).0._State\ is 
                    when \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\BitMask::op_BitwiseOr(BitMask,BitMask).0._Started\ = true) then 
                            \BitMask::op_BitwiseOr(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\BitMask::op_BitwiseOr(BitMask,BitMask).0._Started\ = true) then 
                            \BitMask::op_BitwiseOr(BitMask,BitMask).0._Finished\ <= true;
                        else 
                            \BitMask::op_BitwiseOr(BitMask,BitMask).0._Finished\ <= false;
                            \BitMask::op_BitwiseOr(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_2\ => 
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.left\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0.left.parameter.In\;
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.right\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0.right.parameter.In\;
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.binaryOperationResult.0\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0.left\.\SegmentCount\ /= \BitMask::op_BitwiseOr(BitMask,BitMask).0.right\.\SegmentCount\;
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.flag\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0.binaryOperationResult.0\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_4\ and ends in state \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_5\.
                        --     * The false branch starts in state \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_6\ and ends in state \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_9\.
                        --     * Execution after either branch will continue in the following state: \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_3\.

                        if (\BitMask::op_BitwiseOr(BitMask,BitMask).0.flag\) then 
                            \BitMask::op_BitwiseOr(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_4\;
                        else 
                            \BitMask::op_BitwiseOr(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_3\ => 
                        -- State after the if-else which was started in state \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_2\.
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.return\ <= \BitMask::op_BitwiseOr(BitMask,BitMask).0.result\;
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_4\ => 
                        -- True branch of the if-else started in state \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_2\.
                        -- Initializing record fields to their defaults.
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.result\.\IsNull\ := false;
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.result\.\Size\ := to_unsigned(0, 16);
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.result\.\SegmentCount\ := to_unsigned(0, 16);
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.result\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\ <= \BitMask::op_BitwiseOr(BitMask,BitMask).0.result\;
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\ <= \BitMask::op_BitwiseOr(BitMask,BitMask).0.left\.\Size\;
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\ <= False;
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= true;
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_5\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                        if (\BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ = \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\) then 
                            \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= false;
                            \BitMask::op_BitwiseOr(BitMask,BitMask).0.result\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\;
                            -- Going to the state after the if-else which was started in state \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_2\.
                            if (\BitMask::op_BitwiseOr(BitMask,BitMask).0._State\ = \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_5\) then 
                                \BitMask::op_BitwiseOr(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_3\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_6\ => 
                        -- False branch of the if-else started in state \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_2\.
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.array\ := (others => to_unsigned(0, 32));
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.num\ := to_unsigned(0, 16);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.binaryOperationResult.1\ := resize(signed(\BitMask::op_BitwiseOr(BitMask,BitMask).0.num\), 32) < to_signed(9, 32);
                        if (\BitMask::op_BitwiseOr(BitMask,BitMask).0.binaryOperationResult.1\) then 
                            \BitMask::op_BitwiseOr(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_7\;
                        else 
                            \BitMask::op_BitwiseOr(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_7\ => 
                        -- Repeated state of the while loop which was started in state \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_6\.
                        -- The while loop's condition:
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.binaryOperationResult.2\ := resize(signed(\BitMask::op_BitwiseOr(BitMask,BitMask).0.num\), 32) < to_signed(9, 32);
                        if (\BitMask::op_BitwiseOr(BitMask,BitMask).0.binaryOperationResult.2\) then 
                            \BitMask::op_BitwiseOr(BitMask,BitMask).0.binaryOperationResult.3\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0.left\.\Segments\(to_integer(resize(signed(\BitMask::op_BitwiseOr(BitMask,BitMask).0.num\), 32))) or \BitMask::op_BitwiseOr(BitMask,BitMask).0.right\.\Segments\(to_integer(resize(signed(\BitMask::op_BitwiseOr(BitMask,BitMask).0.num\), 32)));
                            \BitMask::op_BitwiseOr(BitMask,BitMask).0.array\(to_integer(resize(signed(\BitMask::op_BitwiseOr(BitMask,BitMask).0.num\), 32))) := \BitMask::op_BitwiseOr(BitMask,BitMask).0.binaryOperationResult.3\;
                            \BitMask::op_BitwiseOr(BitMask,BitMask).0.binaryOperationResult.4\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0.num\ + to_unsigned(1, 16);
                            \BitMask::op_BitwiseOr(BitMask,BitMask).0.num\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0.binaryOperationResult.4\;
                        else 
                            \BitMask::op_BitwiseOr(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_8\ => 
                        -- State after the while loop which was started in state \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_6\.
                        -- Initializing record fields to their defaults.
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.result\.\IsNull\ := false;
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.result\.\Size\ := to_unsigned(0, 16);
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.result\.\SegmentCount\ := to_unsigned(0, 16);
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.result\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\ <= \BitMask::op_BitwiseOr(BitMask,BitMask).0.result\;
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\ <= \BitMask::op_BitwiseOr(BitMask,BitMask).0.array\;
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= true;
                        \BitMask::op_BitwiseOr(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_9\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_9\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        if (\BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\) then 
                            \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                            \BitMask::op_BitwiseOr(BitMask,BitMask).0.result\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\;
                            \BitMask::op_BitwiseOr(BitMask,BitMask).0.array\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\;
                            -- Going to the state after the if-else which was started in state \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_2\.
                            if (\BitMask::op_BitwiseOr(BitMask,BitMask).0._State\ = \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_9\) then 
                                \BitMask::op_BitwiseOr(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseOr(BitMask,BitMask).0._State_3\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseOr(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseAnd(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 state machine start
    \BitMask::op_BitwiseAnd(BitMask,BitMask).0._StateMachine\: process (\Clock\) 
        Variable \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State\: \BitMask::op_BitwiseAnd(BitMask,BitMask).0._States\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_0\;
        Variable \BitMask::op_BitwiseAnd(BitMask,BitMask).0.left\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_BitwiseAnd(BitMask,BitMask).0.right\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_BitwiseAnd(BitMask,BitMask).0.flag\: boolean := false;
        Variable \BitMask::op_BitwiseAnd(BitMask,BitMask).0.result\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_BitwiseAnd(BitMask,BitMask).0.array\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
        Variable \BitMask::op_BitwiseAnd(BitMask,BitMask).0.num\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_BitwiseAnd(BitMask,BitMask).0.binaryOperationResult.0\: boolean := false;
        Variable \BitMask::op_BitwiseAnd(BitMask,BitMask).0.binaryOperationResult.1\: boolean := false;
        Variable \BitMask::op_BitwiseAnd(BitMask,BitMask).0.binaryOperationResult.2\: boolean := false;
        Variable \BitMask::op_BitwiseAnd(BitMask,BitMask).0.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_BitwiseAnd(BitMask,BitMask).0.binaryOperationResult.4\: unsigned(15 downto 0) := to_unsigned(0, 16);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \BitMask::op_BitwiseAnd(BitMask,BitMask).0._Finished\ <= false;
                \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\ <= false;
                \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= false;
                \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 32));
                \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_0\;
                \BitMask::op_BitwiseAnd(BitMask,BitMask).0.flag\ := false;
                \BitMask::op_BitwiseAnd(BitMask,BitMask).0.array\ := (others => to_unsigned(0, 32));
                \BitMask::op_BitwiseAnd(BitMask,BitMask).0.num\ := to_unsigned(0, 16);
                \BitMask::op_BitwiseAnd(BitMask,BitMask).0.binaryOperationResult.0\ := false;
                \BitMask::op_BitwiseAnd(BitMask,BitMask).0.binaryOperationResult.1\ := false;
                \BitMask::op_BitwiseAnd(BitMask,BitMask).0.binaryOperationResult.2\ := false;
                \BitMask::op_BitwiseAnd(BitMask,BitMask).0.binaryOperationResult.3\ := to_unsigned(0, 32);
                \BitMask::op_BitwiseAnd(BitMask,BitMask).0.binaryOperationResult.4\ := to_unsigned(0, 16);
            else 
                case \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State\ is 
                    when \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\BitMask::op_BitwiseAnd(BitMask,BitMask).0._Started\ = true) then 
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\BitMask::op_BitwiseAnd(BitMask,BitMask).0._Started\ = true) then 
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0._Finished\ <= true;
                        else 
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0._Finished\ <= false;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_2\ => 
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.left\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0.left.parameter.In\;
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.right\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0.right.parameter.In\;
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.binaryOperationResult.0\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0.left\.\SegmentCount\ /= \BitMask::op_BitwiseAnd(BitMask,BitMask).0.right\.\SegmentCount\;
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.flag\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0.binaryOperationResult.0\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_4\ and ends in state \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_5\.
                        --     * The false branch starts in state \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_6\ and ends in state \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_9\.
                        --     * Execution after either branch will continue in the following state: \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_3\.

                        if (\BitMask::op_BitwiseAnd(BitMask,BitMask).0.flag\) then 
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_4\;
                        else 
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_3\ => 
                        -- State after the if-else which was started in state \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_2\.
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.return\ <= \BitMask::op_BitwiseAnd(BitMask,BitMask).0.result\;
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_4\ => 
                        -- True branch of the if-else started in state \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_2\.
                        -- Initializing record fields to their defaults.
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.result\.\IsNull\ := false;
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.result\.\Size\ := to_unsigned(0, 16);
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.result\.\SegmentCount\ := to_unsigned(0, 16);
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.result\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\ <= \BitMask::op_BitwiseAnd(BitMask,BitMask).0.result\;
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\ <= \BitMask::op_BitwiseAnd(BitMask,BitMask).0.left\.\Size\;
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\ <= False;
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= true;
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_5\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                        if (\BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ = \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\) then 
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= false;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.result\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\;
                            -- Going to the state after the if-else which was started in state \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_2\.
                            if (\BitMask::op_BitwiseAnd(BitMask,BitMask).0._State\ = \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_5\) then 
                                \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_3\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_6\ => 
                        -- False branch of the if-else started in state \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_2\.
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.array\ := (others => to_unsigned(0, 32));
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.num\ := to_unsigned(0, 16);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.binaryOperationResult.1\ := resize(signed(\BitMask::op_BitwiseAnd(BitMask,BitMask).0.num\), 32) < to_signed(9, 32);
                        if (\BitMask::op_BitwiseAnd(BitMask,BitMask).0.binaryOperationResult.1\) then 
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_7\;
                        else 
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_7\ => 
                        -- Repeated state of the while loop which was started in state \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_6\.
                        -- The while loop's condition:
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.binaryOperationResult.2\ := resize(signed(\BitMask::op_BitwiseAnd(BitMask,BitMask).0.num\), 32) < to_signed(9, 32);
                        if (\BitMask::op_BitwiseAnd(BitMask,BitMask).0.binaryOperationResult.2\) then 
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.binaryOperationResult.3\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0.left\.\Segments\(to_integer(resize(signed(\BitMask::op_BitwiseAnd(BitMask,BitMask).0.num\), 32))) and \BitMask::op_BitwiseAnd(BitMask,BitMask).0.right\.\Segments\(to_integer(resize(signed(\BitMask::op_BitwiseAnd(BitMask,BitMask).0.num\), 32)));
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.array\(to_integer(resize(signed(\BitMask::op_BitwiseAnd(BitMask,BitMask).0.num\), 32))) := \BitMask::op_BitwiseAnd(BitMask,BitMask).0.binaryOperationResult.3\;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.binaryOperationResult.4\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0.num\ + to_unsigned(1, 16);
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.num\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0.binaryOperationResult.4\;
                        else 
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_8\ => 
                        -- State after the while loop which was started in state \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_6\.
                        -- Initializing record fields to their defaults.
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.result\.\IsNull\ := false;
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.result\.\Size\ := to_unsigned(0, 16);
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.result\.\SegmentCount\ := to_unsigned(0, 16);
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.result\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\ <= \BitMask::op_BitwiseAnd(BitMask,BitMask).0.result\;
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\ <= \BitMask::op_BitwiseAnd(BitMask,BitMask).0.array\;
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= true;
                        \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_9\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_9\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        if (\BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\) then 
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.result\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.array\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\;
                            -- Going to the state after the if-else which was started in state \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_2\.
                            if (\BitMask::op_BitwiseAnd(BitMask,BitMask).0._State\ = \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_9\) then 
                                \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State\ := \BitMask::op_BitwiseAnd(BitMask,BitMask).0._State_3\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseAnd(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_RightShift(Lombiq.Unum.BitMask,System.Int32).0 state machine start
    \BitMask::op_RightShift(BitMask,Int32).0._StateMachine\: process (\Clock\) 
        Variable \BitMask::op_RightShift(BitMask,Int32).0._State\: \BitMask::op_RightShift(BitMask,Int32).0._States\ := \BitMask::op_RightShift(BitMask,Int32).0._State_0\;
        Variable \BitMask::op_RightShift(BitMask,Int32).0.left\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_RightShift(BitMask,Int32).0.right\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_RightShift(BitMask,Int32).0.flag\: boolean := false;
        Variable \BitMask::op_RightShift(BitMask,Int32).0.result\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_RightShift(BitMask,Int32).0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_RightShift(BitMask,Int32).0.array\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
        Variable \BitMask::op_RightShift(BitMask,Int32).0.num2\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_RightShift(BitMask,Int32).0.flag2\: boolean := false;
        Variable \BitMask::op_RightShift(BitMask,Int32).0.num3\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_RightShift(BitMask,Int32).0.num4\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_RightShift(BitMask,Int32).0.flag3\: boolean := false;
        Variable \BitMask::op_RightShift(BitMask,Int32).0.flag4\: boolean := false;
        Variable \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.0\: boolean := false;
        Variable \BitMask::op_RightShift(BitMask,Int32).0.return.0\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.1\: boolean := false;
        Variable \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.2\: boolean := false;
        Variable \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.3\: boolean := false;
        Variable \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.4\: boolean := false;
        Variable \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.5\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.6\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_RightShift(BitMask,Int32).0.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.7\: boolean := false;
        Variable \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.8\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.9\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.10\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.11\: unsigned(15 downto 0) := to_unsigned(0, 16);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \BitMask::op_RightShift(BitMask,Int32).0._Finished\ <= false;
                \BitMask::op_RightShift(BitMask,Int32).0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\ <= to_signed(0, 32);
                \BitMask::op_RightShift(BitMask,Int32).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= false;
                \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 32));
                \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                \BitMask::op_RightShift(BitMask,Int32).0._State\ := \BitMask::op_RightShift(BitMask,Int32).0._State_0\;
                \BitMask::op_RightShift(BitMask,Int32).0.right\ := to_signed(0, 32);
                \BitMask::op_RightShift(BitMask,Int32).0.flag\ := false;
                \BitMask::op_RightShift(BitMask,Int32).0.num\ := to_unsigned(0, 32);
                \BitMask::op_RightShift(BitMask,Int32).0.array\ := (others => to_unsigned(0, 32));
                \BitMask::op_RightShift(BitMask,Int32).0.num2\ := to_unsigned(0, 16);
                \BitMask::op_RightShift(BitMask,Int32).0.flag2\ := false;
                \BitMask::op_RightShift(BitMask,Int32).0.num3\ := to_unsigned(0, 16);
                \BitMask::op_RightShift(BitMask,Int32).0.num4\ := to_unsigned(0, 16);
                \BitMask::op_RightShift(BitMask,Int32).0.flag3\ := false;
                \BitMask::op_RightShift(BitMask,Int32).0.flag4\ := false;
                \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.0\ := false;
                \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.1\ := false;
                \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.2\ := false;
                \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.3\ := false;
                \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.4\ := false;
                \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.5\ := to_unsigned(0, 16);
                \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.6\ := to_unsigned(0, 32);
                \BitMask::op_RightShift(BitMask,Int32).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.7\ := false;
                \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.8\ := to_unsigned(0, 32);
                \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.9\ := to_unsigned(0, 32);
                \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.10\ := to_unsigned(0, 16);
                \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.11\ := to_unsigned(0, 16);
            else 
                case \BitMask::op_RightShift(BitMask,Int32).0._State\ is 
                    when \BitMask::op_RightShift(BitMask,Int32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\BitMask::op_RightShift(BitMask,Int32).0._Started\ = true) then 
                            \BitMask::op_RightShift(BitMask,Int32).0._State\ := \BitMask::op_RightShift(BitMask,Int32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_RightShift(BitMask,Int32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\BitMask::op_RightShift(BitMask,Int32).0._Started\ = true) then 
                            \BitMask::op_RightShift(BitMask,Int32).0._Finished\ <= true;
                        else 
                            \BitMask::op_RightShift(BitMask,Int32).0._Finished\ <= false;
                            \BitMask::op_RightShift(BitMask,Int32).0._State\ := \BitMask::op_RightShift(BitMask,Int32).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_RightShift(BitMask,Int32).0._State_2\ => 
                        \BitMask::op_RightShift(BitMask,Int32).0.left\ := \BitMask::op_RightShift(BitMask,Int32).0.left.parameter.In\;
                        \BitMask::op_RightShift(BitMask,Int32).0.right\ := \BitMask::op_RightShift(BitMask,Int32).0.right.parameter.In\;
                        \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.0\ := \BitMask::op_RightShift(BitMask,Int32).0.right\ < to_signed(0, 32);
                        \BitMask::op_RightShift(BitMask,Int32).0.flag\ := \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.0\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::op_RightShift(BitMask,Int32).0._State_4\ and ends in state \BitMask::op_RightShift(BitMask,Int32).0._State_5\.
                        --     * The false branch starts in state \BitMask::op_RightShift(BitMask,Int32).0._State_6\ and ends in state \BitMask::op_RightShift(BitMask,Int32).0._State_15\.
                        --     * Execution after either branch will continue in the following state: \BitMask::op_RightShift(BitMask,Int32).0._State_3\.

                        if (\BitMask::op_RightShift(BitMask,Int32).0.flag\) then 
                            \BitMask::op_RightShift(BitMask,Int32).0._State\ := \BitMask::op_RightShift(BitMask,Int32).0._State_4\;
                        else 
                            \BitMask::op_RightShift(BitMask,Int32).0._State\ := \BitMask::op_RightShift(BitMask,Int32).0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_RightShift(BitMask,Int32).0._State_3\ => 
                        -- State after the if-else which was started in state \BitMask::op_RightShift(BitMask,Int32).0._State_2\.
                        \BitMask::op_RightShift(BitMask,Int32).0.return\ <= \BitMask::op_RightShift(BitMask,Int32).0.result\;
                        \BitMask::op_RightShift(BitMask,Int32).0._State\ := \BitMask::op_RightShift(BitMask,Int32).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_RightShift(BitMask,Int32).0._State_4\ => 
                        -- True branch of the if-else started in state \BitMask::op_RightShift(BitMask,Int32).0._State_2\.
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                        \BitMask::op_RightShift(BitMask,Int32).0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\ <= \BitMask::op_RightShift(BitMask,Int32).0.left\;
                        \BitMask::op_RightShift(BitMask,Int32).0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\ <= -\BitMask::op_RightShift(BitMask,Int32).0.right\;
                        \BitMask::op_RightShift(BitMask,Int32).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= true;
                        \BitMask::op_RightShift(BitMask,Int32).0._State\ := \BitMask::op_RightShift(BitMask,Int32).0._State_5\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_RightShift(BitMask,Int32).0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                        if (\BitMask::op_RightShift(BitMask,Int32).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ = \BitMask::op_RightShift(BitMask,Int32).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\) then 
                            \BitMask::op_RightShift(BitMask,Int32).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= false;
                            \BitMask::op_RightShift(BitMask,Int32).0.return.0\ := \BitMask::op_RightShift(BitMask,Int32).0.BitMask::op_LeftShift(BitMask,Int32).return.0\;
                            \BitMask::op_RightShift(BitMask,Int32).0.result\ := \BitMask::op_RightShift(BitMask,Int32).0.return.0\;
                            -- Going to the state after the if-else which was started in state \BitMask::op_RightShift(BitMask,Int32).0._State_2\.
                            if (\BitMask::op_RightShift(BitMask,Int32).0._State\ = \BitMask::op_RightShift(BitMask,Int32).0._State_5\) then 
                                \BitMask::op_RightShift(BitMask,Int32).0._State\ := \BitMask::op_RightShift(BitMask,Int32).0._State_3\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_RightShift(BitMask,Int32).0._State_6\ => 
                        -- False branch of the if-else started in state \BitMask::op_RightShift(BitMask,Int32).0._State_2\.
                        -- Since the integer literal 2147483648 was out of the VHDL integer range it was substituted with a binary literal (10000000000000000000000000000000).
                        \BitMask::op_RightShift(BitMask,Int32).0.num\ := "10000000000000000000000000000000";
                        \BitMask::op_RightShift(BitMask,Int32).0.array\ := (others => to_unsigned(0, 32));
                        \BitMask::op_RightShift(BitMask,Int32).0.array\ := \BitMask::op_RightShift(BitMask,Int32).0.left\.\Segments\(0 to 8);
                        \BitMask::op_RightShift(BitMask,Int32).0.num2\ := to_unsigned(0, 16);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.1\ := resize(signed(\BitMask::op_RightShift(BitMask,Int32).0.num2\), 32) < \BitMask::op_RightShift(BitMask,Int32).0.right\;
                        if (\BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.1\) then 
                            \BitMask::op_RightShift(BitMask,Int32).0._State\ := \BitMask::op_RightShift(BitMask,Int32).0._State_7\;
                        else 
                            \BitMask::op_RightShift(BitMask,Int32).0._State\ := \BitMask::op_RightShift(BitMask,Int32).0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_RightShift(BitMask,Int32).0._State_7\ => 
                        -- Repeated state of the while loop which was started in state \BitMask::op_RightShift(BitMask,Int32).0._State_6\.
                        -- The while loop's condition:
                        \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.2\ := resize(signed(\BitMask::op_RightShift(BitMask,Int32).0.num2\), 32) < \BitMask::op_RightShift(BitMask,Int32).0.right\;
                        if (\BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.2\) then 
                            \BitMask::op_RightShift(BitMask,Int32).0.flag2\ := False;
                            \BitMask::op_RightShift(BitMask,Int32).0.num3\ := to_unsigned(1, 16);
                            -- Starting a while loop.
                            -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                            \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.3\ := resize(signed(\BitMask::op_RightShift(BitMask,Int32).0.num3\), 32) <= to_signed(9, 32);
                            if (\BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.3\) then 
                                \BitMask::op_RightShift(BitMask,Int32).0._State\ := \BitMask::op_RightShift(BitMask,Int32).0._State_9\;
                            else 
                                \BitMask::op_RightShift(BitMask,Int32).0._State\ := \BitMask::op_RightShift(BitMask,Int32).0._State_10\;
                            end if;
                        else 
                            \BitMask::op_RightShift(BitMask,Int32).0._State\ := \BitMask::op_RightShift(BitMask,Int32).0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \BitMask::op_RightShift(BitMask,Int32).0._State_8\ => 
                        -- State after the while loop which was started in state \BitMask::op_RightShift(BitMask,Int32).0._State_6\.
                        -- Initializing record fields to their defaults.
                        \BitMask::op_RightShift(BitMask,Int32).0.result\.\IsNull\ := false;
                        \BitMask::op_RightShift(BitMask,Int32).0.result\.\Size\ := to_unsigned(0, 16);
                        \BitMask::op_RightShift(BitMask,Int32).0.result\.\SegmentCount\ := to_unsigned(0, 16);
                        \BitMask::op_RightShift(BitMask,Int32).0.result\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\ <= \BitMask::op_RightShift(BitMask,Int32).0.result\;
                        \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\ <= \BitMask::op_RightShift(BitMask,Int32).0.array\;
                        \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                        \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= true;
                        \BitMask::op_RightShift(BitMask,Int32).0._State\ := \BitMask::op_RightShift(BitMask,Int32).0._State_15\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_RightShift(BitMask,Int32).0._State_9\ => 
                        -- Repeated state of the while loop which was started in state \BitMask::op_RightShift(BitMask,Int32).0._State_7\.
                        -- The while loop's condition:
                        \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.4\ := resize(signed(\BitMask::op_RightShift(BitMask,Int32).0.num3\), 32) <= to_signed(9, 32);
                        if (\BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.4\) then 
                            \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.5\ := resize(unsigned(to_signed(9, 32) - resize(signed(\BitMask::op_RightShift(BitMask,Int32).0.num3\), 32)), 16);
                            \BitMask::op_RightShift(BitMask,Int32).0.num4\ := (\BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.5\);
                            \BitMask::op_RightShift(BitMask,Int32).0._State\ := \BitMask::op_RightShift(BitMask,Int32).0._State_11\;
                        else 
                            \BitMask::op_RightShift(BitMask,Int32).0._State\ := \BitMask::op_RightShift(BitMask,Int32).0._State_10\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \BitMask::op_RightShift(BitMask,Int32).0._State_10\ => 
                        -- State after the while loop which was started in state \BitMask::op_RightShift(BitMask,Int32).0._State_7\.
                        \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.11\ := \BitMask::op_RightShift(BitMask,Int32).0.num2\ + to_unsigned(1, 16);
                        \BitMask::op_RightShift(BitMask,Int32).0.num2\ := \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.11\;
                        -- Returning to the repeated state of the while loop which was started in state \BitMask::op_RightShift(BitMask,Int32).0._State_6\ if the loop wasn't exited with a state change.
                        if (\BitMask::op_RightShift(BitMask,Int32).0._State\ = \BitMask::op_RightShift(BitMask,Int32).0._State_10\) then 
                            \BitMask::op_RightShift(BitMask,Int32).0._State\ := \BitMask::op_RightShift(BitMask,Int32).0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_RightShift(BitMask,Int32).0._State_11\ => 
                        -- Waiting for the result to appear in \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.6\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\BitMask::op_RightShift(BitMask,Int32).0.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \BitMask::op_RightShift(BitMask,Int32).0._State\ := \BitMask::op_RightShift(BitMask,Int32).0._State_12\;
                            \BitMask::op_RightShift(BitMask,Int32).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \BitMask::op_RightShift(BitMask,Int32).0.clockCyclesWaitedForBinaryOperationResult.0\ := \BitMask::op_RightShift(BitMask,Int32).0.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.6\ := \BitMask::op_RightShift(BitMask,Int32).0.array\(to_integer(resize(signed(\BitMask::op_RightShift(BitMask,Int32).0.num4\), 32))) mod to_unsigned(2, 32);
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \BitMask::op_RightShift(BitMask,Int32).0._State_12\ => 
                        \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.7\ := \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.6\ = to_unsigned(1, 32);
                        \BitMask::op_RightShift(BitMask,Int32).0.flag3\ := \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.7\;
                        \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.8\ := shift_right(\BitMask::op_RightShift(BitMask,Int32).0.array\(to_integer(resize(signed(\BitMask::op_RightShift(BitMask,Int32).0.num4\), 32))), to_integer(to_signed(1, 32)));
                        \BitMask::op_RightShift(BitMask,Int32).0.array\(to_integer(resize(signed(\BitMask::op_RightShift(BitMask,Int32).0.num4\), 32))) := \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.8\;
                        \BitMask::op_RightShift(BitMask,Int32).0.flag4\ := \BitMask::op_RightShift(BitMask,Int32).0.flag2\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::op_RightShift(BitMask,Int32).0._State_14\ and ends in state \BitMask::op_RightShift(BitMask,Int32).0._State_14\.
                        --     * Execution after either branch will continue in the following state: \BitMask::op_RightShift(BitMask,Int32).0._State_13\.

                        if (\BitMask::op_RightShift(BitMask,Int32).0.flag4\) then 
                            \BitMask::op_RightShift(BitMask,Int32).0._State\ := \BitMask::op_RightShift(BitMask,Int32).0._State_14\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \BitMask::op_RightShift(BitMask,Int32).0._State\ := \BitMask::op_RightShift(BitMask,Int32).0._State_13\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \BitMask::op_RightShift(BitMask,Int32).0._State_13\ => 
                        -- State after the if-else which was started in state \BitMask::op_RightShift(BitMask,Int32).0._State_12\.
                        \BitMask::op_RightShift(BitMask,Int32).0.flag2\ := \BitMask::op_RightShift(BitMask,Int32).0.flag3\;
                        \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.10\ := \BitMask::op_RightShift(BitMask,Int32).0.num3\ + to_unsigned(1, 16);
                        \BitMask::op_RightShift(BitMask,Int32).0.num3\ := \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.10\;
                        -- Returning to the repeated state of the while loop which was started in state \BitMask::op_RightShift(BitMask,Int32).0._State_7\ if the loop wasn't exited with a state change.
                        if (\BitMask::op_RightShift(BitMask,Int32).0._State\ = \BitMask::op_RightShift(BitMask,Int32).0._State_13\) then 
                            \BitMask::op_RightShift(BitMask,Int32).0._State\ := \BitMask::op_RightShift(BitMask,Int32).0._State_9\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_RightShift(BitMask,Int32).0._State_14\ => 
                        -- True branch of the if-else started in state \BitMask::op_RightShift(BitMask,Int32).0._State_12\.
                        \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.9\ := \BitMask::op_RightShift(BitMask,Int32).0.array\(to_integer(resize(signed(\BitMask::op_RightShift(BitMask,Int32).0.num4\), 32))) or \BitMask::op_RightShift(BitMask,Int32).0.num\;
                        \BitMask::op_RightShift(BitMask,Int32).0.array\(to_integer(resize(signed(\BitMask::op_RightShift(BitMask,Int32).0.num4\), 32))) := \BitMask::op_RightShift(BitMask,Int32).0.binaryOperationResult.9\;
                        -- Going to the state after the if-else which was started in state \BitMask::op_RightShift(BitMask,Int32).0._State_12\.
                        if (\BitMask::op_RightShift(BitMask,Int32).0._State\ = \BitMask::op_RightShift(BitMask,Int32).0._State_14\) then 
                            \BitMask::op_RightShift(BitMask,Int32).0._State\ := \BitMask::op_RightShift(BitMask,Int32).0._State_13\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_RightShift(BitMask,Int32).0._State_15\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        if (\BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\) then 
                            \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                            \BitMask::op_RightShift(BitMask,Int32).0.result\ := \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\;
                            \BitMask::op_RightShift(BitMask,Int32).0.array\ := \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\;
                            -- Going to the state after the if-else which was started in state \BitMask::op_RightShift(BitMask,Int32).0._State_2\.
                            if (\BitMask::op_RightShift(BitMask,Int32).0._State\ = \BitMask::op_RightShift(BitMask,Int32).0._State_15\) then 
                                \BitMask::op_RightShift(BitMask,Int32).0._State\ := \BitMask::op_RightShift(BitMask,Int32).0._State_3\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_RightShift(Lombiq.Unum.BitMask,System.Int32).0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32).0 state machine start
    \BitMask::op_LeftShift(BitMask,Int32).0._StateMachine\: process (\Clock\) 
        Variable \BitMask::op_LeftShift(BitMask,Int32).0._State\: \BitMask::op_LeftShift(BitMask,Int32).0._States\ := \BitMask::op_LeftShift(BitMask,Int32).0._State_0\;
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.left\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.right\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.flag\: boolean := false;
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.result\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.num2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.array\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.num3\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.flag2\: boolean := false;
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.num4\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.flag3\: boolean := false;
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.flag4\: boolean := false;
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.0\: boolean := false;
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.return.0\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.1\: boolean := false;
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.2\: boolean := false;
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.3\: boolean := false;
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.4\: boolean := false;
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.5\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.6\: boolean := false;
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.7\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.8\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.9\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.10\: unsigned(15 downto 0) := to_unsigned(0, 16);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \BitMask::op_LeftShift(BitMask,Int32).0._Finished\ <= false;
                \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::op_RightShift(BitMask,Int32).right.parameter.Out.0\ <= to_signed(0, 32);
                \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ <= false;
                \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 32));
                \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                \BitMask::op_LeftShift(BitMask,Int32).0._State\ := \BitMask::op_LeftShift(BitMask,Int32).0._State_0\;
                \BitMask::op_LeftShift(BitMask,Int32).0.right\ := to_signed(0, 32);
                \BitMask::op_LeftShift(BitMask,Int32).0.flag\ := false;
                \BitMask::op_LeftShift(BitMask,Int32).0.num\ := to_unsigned(0, 32);
                \BitMask::op_LeftShift(BitMask,Int32).0.num2\ := to_unsigned(0, 32);
                \BitMask::op_LeftShift(BitMask,Int32).0.array\ := (others => to_unsigned(0, 32));
                \BitMask::op_LeftShift(BitMask,Int32).0.num3\ := to_unsigned(0, 16);
                \BitMask::op_LeftShift(BitMask,Int32).0.flag2\ := false;
                \BitMask::op_LeftShift(BitMask,Int32).0.num4\ := to_unsigned(0, 16);
                \BitMask::op_LeftShift(BitMask,Int32).0.flag3\ := false;
                \BitMask::op_LeftShift(BitMask,Int32).0.flag4\ := false;
                \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.0\ := false;
                \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.1\ := false;
                \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.2\ := false;
                \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.3\ := false;
                \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.4\ := false;
                \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.5\ := to_unsigned(0, 32);
                \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.6\ := false;
                \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.7\ := to_unsigned(0, 32);
                \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.8\ := to_unsigned(0, 32);
                \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.9\ := to_unsigned(0, 16);
                \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.10\ := to_unsigned(0, 16);
            else 
                case \BitMask::op_LeftShift(BitMask,Int32).0._State\ is 
                    when \BitMask::op_LeftShift(BitMask,Int32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\BitMask::op_LeftShift(BitMask,Int32).0._Started\ = true) then 
                            \BitMask::op_LeftShift(BitMask,Int32).0._State\ := \BitMask::op_LeftShift(BitMask,Int32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_LeftShift(BitMask,Int32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\BitMask::op_LeftShift(BitMask,Int32).0._Started\ = true) then 
                            \BitMask::op_LeftShift(BitMask,Int32).0._Finished\ <= true;
                        else 
                            \BitMask::op_LeftShift(BitMask,Int32).0._Finished\ <= false;
                            \BitMask::op_LeftShift(BitMask,Int32).0._State\ := \BitMask::op_LeftShift(BitMask,Int32).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_LeftShift(BitMask,Int32).0._State_2\ => 
                        \BitMask::op_LeftShift(BitMask,Int32).0.left\ := \BitMask::op_LeftShift(BitMask,Int32).0.left.parameter.In\;
                        \BitMask::op_LeftShift(BitMask,Int32).0.right\ := \BitMask::op_LeftShift(BitMask,Int32).0.right.parameter.In\;
                        \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.0\ := \BitMask::op_LeftShift(BitMask,Int32).0.right\ < to_signed(0, 32);
                        \BitMask::op_LeftShift(BitMask,Int32).0.flag\ := \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.0\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::op_LeftShift(BitMask,Int32).0._State_4\ and ends in state \BitMask::op_LeftShift(BitMask,Int32).0._State_5\.
                        --     * The false branch starts in state \BitMask::op_LeftShift(BitMask,Int32).0._State_6\ and ends in state \BitMask::op_LeftShift(BitMask,Int32).0._State_13\.
                        --     * Execution after either branch will continue in the following state: \BitMask::op_LeftShift(BitMask,Int32).0._State_3\.

                        if (\BitMask::op_LeftShift(BitMask,Int32).0.flag\) then 
                            \BitMask::op_LeftShift(BitMask,Int32).0._State\ := \BitMask::op_LeftShift(BitMask,Int32).0._State_4\;
                        else 
                            \BitMask::op_LeftShift(BitMask,Int32).0._State\ := \BitMask::op_LeftShift(BitMask,Int32).0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_LeftShift(BitMask,Int32).0._State_3\ => 
                        -- State after the if-else which was started in state \BitMask::op_LeftShift(BitMask,Int32).0._State_2\.
                        \BitMask::op_LeftShift(BitMask,Int32).0.return\ <= \BitMask::op_LeftShift(BitMask,Int32).0.result\;
                        \BitMask::op_LeftShift(BitMask,Int32).0._State\ := \BitMask::op_LeftShift(BitMask,Int32).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_LeftShift(BitMask,Int32).0._State_4\ => 
                        -- True branch of the if-else started in state \BitMask::op_LeftShift(BitMask,Int32).0._State_2\.
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_RightShift(Lombiq.Unum.BitMask,System.Int32)
                        \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::op_RightShift(BitMask,Int32).left.parameter.Out.0\ <= \BitMask::op_LeftShift(BitMask,Int32).0.left\;
                        \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::op_RightShift(BitMask,Int32).right.parameter.Out.0\ <= -\BitMask::op_LeftShift(BitMask,Int32).0.right\;
                        \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ <= true;
                        \BitMask::op_LeftShift(BitMask,Int32).0._State\ := \BitMask::op_LeftShift(BitMask,Int32).0._State_5\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_LeftShift(BitMask,Int32).0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_RightShift(Lombiq.Unum.BitMask,System.Int32)
                        if (\BitMask::op_LeftShift(BitMask,Int32).0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ = \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\) then 
                            \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ <= false;
                            \BitMask::op_LeftShift(BitMask,Int32).0.return.0\ := \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::op_RightShift(BitMask,Int32).return.0\;
                            \BitMask::op_LeftShift(BitMask,Int32).0.result\ := \BitMask::op_LeftShift(BitMask,Int32).0.return.0\;
                            -- Going to the state after the if-else which was started in state \BitMask::op_LeftShift(BitMask,Int32).0._State_2\.
                            if (\BitMask::op_LeftShift(BitMask,Int32).0._State\ = \BitMask::op_LeftShift(BitMask,Int32).0._State_5\) then 
                                \BitMask::op_LeftShift(BitMask,Int32).0._State\ := \BitMask::op_LeftShift(BitMask,Int32).0._State_3\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_LeftShift(BitMask,Int32).0._State_6\ => 
                        -- False branch of the if-else started in state \BitMask::op_LeftShift(BitMask,Int32).0._State_2\.
                        -- Since the integer literal 2147483648 was out of the VHDL integer range it was substituted with a binary literal (10000000000000000000000000000000).
                        \BitMask::op_LeftShift(BitMask,Int32).0.num\ := "10000000000000000000000000000000";
                        \BitMask::op_LeftShift(BitMask,Int32).0.num2\ := to_unsigned(1, 32);
                        \BitMask::op_LeftShift(BitMask,Int32).0.array\ := (others => to_unsigned(0, 32));
                        \BitMask::op_LeftShift(BitMask,Int32).0.array\ := \BitMask::op_LeftShift(BitMask,Int32).0.left\.\Segments\(0 to 8);
                        \BitMask::op_LeftShift(BitMask,Int32).0.num3\ := to_unsigned(0, 16);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.1\ := resize(signed(\BitMask::op_LeftShift(BitMask,Int32).0.num3\), 32) < \BitMask::op_LeftShift(BitMask,Int32).0.right\;
                        if (\BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.1\) then 
                            \BitMask::op_LeftShift(BitMask,Int32).0._State\ := \BitMask::op_LeftShift(BitMask,Int32).0._State_7\;
                        else 
                            \BitMask::op_LeftShift(BitMask,Int32).0._State\ := \BitMask::op_LeftShift(BitMask,Int32).0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_LeftShift(BitMask,Int32).0._State_7\ => 
                        -- Repeated state of the while loop which was started in state \BitMask::op_LeftShift(BitMask,Int32).0._State_6\.
                        -- The while loop's condition:
                        \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.2\ := resize(signed(\BitMask::op_LeftShift(BitMask,Int32).0.num3\), 32) < \BitMask::op_LeftShift(BitMask,Int32).0.right\;
                        if (\BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.2\) then 
                            \BitMask::op_LeftShift(BitMask,Int32).0.flag2\ := False;
                            \BitMask::op_LeftShift(BitMask,Int32).0.num4\ := to_unsigned(0, 16);
                            -- Starting a while loop.
                            -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                            \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.3\ := resize(signed(\BitMask::op_LeftShift(BitMask,Int32).0.num4\), 32) < to_signed(9, 32);
                            if (\BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.3\) then 
                                \BitMask::op_LeftShift(BitMask,Int32).0._State\ := \BitMask::op_LeftShift(BitMask,Int32).0._State_9\;
                            else 
                                \BitMask::op_LeftShift(BitMask,Int32).0._State\ := \BitMask::op_LeftShift(BitMask,Int32).0._State_10\;
                            end if;
                        else 
                            \BitMask::op_LeftShift(BitMask,Int32).0._State\ := \BitMask::op_LeftShift(BitMask,Int32).0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \BitMask::op_LeftShift(BitMask,Int32).0._State_8\ => 
                        -- State after the while loop which was started in state \BitMask::op_LeftShift(BitMask,Int32).0._State_6\.
                        -- Initializing record fields to their defaults.
                        \BitMask::op_LeftShift(BitMask,Int32).0.result\.\IsNull\ := false;
                        \BitMask::op_LeftShift(BitMask,Int32).0.result\.\Size\ := to_unsigned(0, 16);
                        \BitMask::op_LeftShift(BitMask,Int32).0.result\.\SegmentCount\ := to_unsigned(0, 16);
                        \BitMask::op_LeftShift(BitMask,Int32).0.result\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\ <= \BitMask::op_LeftShift(BitMask,Int32).0.result\;
                        \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\ <= \BitMask::op_LeftShift(BitMask,Int32).0.array\;
                        \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                        \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= true;
                        \BitMask::op_LeftShift(BitMask,Int32).0._State\ := \BitMask::op_LeftShift(BitMask,Int32).0._State_13\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::op_LeftShift(BitMask,Int32).0._State_9\ => 
                        -- Repeated state of the while loop which was started in state \BitMask::op_LeftShift(BitMask,Int32).0._State_7\.
                        -- The while loop's condition:
                        \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.4\ := resize(signed(\BitMask::op_LeftShift(BitMask,Int32).0.num4\), 32) < to_signed(9, 32);
                        if (\BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.4\) then 
                            \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.5\ := \BitMask::op_LeftShift(BitMask,Int32).0.array\(to_integer(resize(signed(\BitMask::op_LeftShift(BitMask,Int32).0.num4\), 32))) and \BitMask::op_LeftShift(BitMask,Int32).0.num\;
                            \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.6\ := \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.5\ = \BitMask::op_LeftShift(BitMask,Int32).0.num\;
                            \BitMask::op_LeftShift(BitMask,Int32).0.flag3\ := \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.6\;
                            \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.7\ := shift_left(\BitMask::op_LeftShift(BitMask,Int32).0.array\(to_integer(resize(signed(\BitMask::op_LeftShift(BitMask,Int32).0.num4\), 32))), to_integer(to_signed(1, 32)));
                            \BitMask::op_LeftShift(BitMask,Int32).0.array\(to_integer(resize(signed(\BitMask::op_LeftShift(BitMask,Int32).0.num4\), 32))) := \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.7\;
                            \BitMask::op_LeftShift(BitMask,Int32).0.flag4\ := \BitMask::op_LeftShift(BitMask,Int32).0.flag2\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \BitMask::op_LeftShift(BitMask,Int32).0._State_12\ and ends in state \BitMask::op_LeftShift(BitMask,Int32).0._State_12\.
                            --     * Execution after either branch will continue in the following state: \BitMask::op_LeftShift(BitMask,Int32).0._State_11\.

                            if (\BitMask::op_LeftShift(BitMask,Int32).0.flag4\) then 
                                \BitMask::op_LeftShift(BitMask,Int32).0._State\ := \BitMask::op_LeftShift(BitMask,Int32).0._State_12\;
                            else 
                                -- There was no false branch, so going directly to the state after the if-else.
                                \BitMask::op_LeftShift(BitMask,Int32).0._State\ := \BitMask::op_LeftShift(BitMask,Int32).0._State_11\;
                            end if;
                        else 
                            \BitMask::op_LeftShift(BitMask,Int32).0._State\ := \BitMask::op_LeftShift(BitMask,Int32).0._State_10\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.4
                    when \BitMask::op_LeftShift(BitMask,Int32).0._State_10\ => 
                        -- State after the while loop which was started in state \BitMask::op_LeftShift(BitMask,Int32).0._State_7\.
                        \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.10\ := \BitMask::op_LeftShift(BitMask,Int32).0.num3\ + to_unsigned(1, 16);
                        \BitMask::op_LeftShift(BitMask,Int32).0.num3\ := \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.10\;
                        -- Returning to the repeated state of the while loop which was started in state \BitMask::op_LeftShift(BitMask,Int32).0._State_6\ if the loop wasn't exited with a state change.
                        if (\BitMask::op_LeftShift(BitMask,Int32).0._State\ = \BitMask::op_LeftShift(BitMask,Int32).0._State_10\) then 
                            \BitMask::op_LeftShift(BitMask,Int32).0._State\ := \BitMask::op_LeftShift(BitMask,Int32).0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_LeftShift(BitMask,Int32).0._State_11\ => 
                        -- State after the if-else which was started in state \BitMask::op_LeftShift(BitMask,Int32).0._State_9\.
                        \BitMask::op_LeftShift(BitMask,Int32).0.flag2\ := \BitMask::op_LeftShift(BitMask,Int32).0.flag3\;
                        \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.9\ := \BitMask::op_LeftShift(BitMask,Int32).0.num4\ + to_unsigned(1, 16);
                        \BitMask::op_LeftShift(BitMask,Int32).0.num4\ := \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.9\;
                        -- Returning to the repeated state of the while loop which was started in state \BitMask::op_LeftShift(BitMask,Int32).0._State_7\ if the loop wasn't exited with a state change.
                        if (\BitMask::op_LeftShift(BitMask,Int32).0._State\ = \BitMask::op_LeftShift(BitMask,Int32).0._State_11\) then 
                            \BitMask::op_LeftShift(BitMask,Int32).0._State\ := \BitMask::op_LeftShift(BitMask,Int32).0._State_9\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_LeftShift(BitMask,Int32).0._State_12\ => 
                        -- True branch of the if-else started in state \BitMask::op_LeftShift(BitMask,Int32).0._State_9\.
                        \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.8\ := \BitMask::op_LeftShift(BitMask,Int32).0.array\(to_integer(resize(signed(\BitMask::op_LeftShift(BitMask,Int32).0.num4\), 32))) or \BitMask::op_LeftShift(BitMask,Int32).0.num2\;
                        \BitMask::op_LeftShift(BitMask,Int32).0.array\(to_integer(resize(signed(\BitMask::op_LeftShift(BitMask,Int32).0.num4\), 32))) := \BitMask::op_LeftShift(BitMask,Int32).0.binaryOperationResult.8\;
                        -- Going to the state after the if-else which was started in state \BitMask::op_LeftShift(BitMask,Int32).0._State_9\.
                        if (\BitMask::op_LeftShift(BitMask,Int32).0._State\ = \BitMask::op_LeftShift(BitMask,Int32).0._State_12\) then 
                            \BitMask::op_LeftShift(BitMask,Int32).0._State\ := \BitMask::op_LeftShift(BitMask,Int32).0._State_11\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::op_LeftShift(BitMask,Int32).0._State_13\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        if (\BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\) then 
                            \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                            \BitMask::op_LeftShift(BitMask,Int32).0.result\ := \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\;
                            \BitMask::op_LeftShift(BitMask,Int32).0.array\ := \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\;
                            -- Going to the state after the if-else which was started in state \BitMask::op_LeftShift(BitMask,Int32).0._State_2\.
                            if (\BitMask::op_LeftShift(BitMask,Int32).0._State\ = \BitMask::op_LeftShift(BitMask,Int32).0._State_13\) then 
                                \BitMask::op_LeftShift(BitMask,Int32).0._State\ := \BitMask::op_LeftShift(BitMask,Int32).0._State_3\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32).0 state machine end


    -- System.UInt16 Lombiq.Unum.BitMask::GetMostSignificantOnePosition().0 state machine start
    \BitMask::GetMostSignificantOnePosition().0._StateMachine\: process (\Clock\) 
        Variable \BitMask::GetMostSignificantOnePosition().0._State\: \BitMask::GetMostSignificantOnePosition().0._States\ := \BitMask::GetMostSignificantOnePosition().0._State_0\;
        Variable \BitMask::GetMostSignificantOnePosition().0.this\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::GetMostSignificantOnePosition().0.num\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::GetMostSignificantOnePosition().0.num2\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::GetMostSignificantOnePosition().0.num3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::GetMostSignificantOnePosition().0.flag\: boolean := false;
        Variable \BitMask::GetMostSignificantOnePosition().0.result\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.0\: boolean := false;
        Variable \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.1\: boolean := false;
        Variable \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.3\: boolean := false;
        Variable \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.4\: boolean := false;
        Variable \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.5\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.6\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.7\: boolean := false;
        Variable \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.8\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.9\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.10\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.11\: unsigned(15 downto 0) := to_unsigned(0, 16);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \BitMask::GetMostSignificantOnePosition().0._Finished\ <= false;
                \BitMask::GetMostSignificantOnePosition().0.return\ <= to_unsigned(0, 16);
                \BitMask::GetMostSignificantOnePosition().0._State\ := \BitMask::GetMostSignificantOnePosition().0._State_0\;
                \BitMask::GetMostSignificantOnePosition().0.num\ := to_unsigned(0, 16);
                \BitMask::GetMostSignificantOnePosition().0.num2\ := to_unsigned(0, 16);
                \BitMask::GetMostSignificantOnePosition().0.num3\ := to_unsigned(0, 32);
                \BitMask::GetMostSignificantOnePosition().0.flag\ := false;
                \BitMask::GetMostSignificantOnePosition().0.result\ := to_unsigned(0, 16);
                \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.0\ := false;
                \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.1\ := false;
                \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.2\ := to_signed(0, 32);
                \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.3\ := false;
                \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.4\ := false;
                \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.5\ := to_unsigned(0, 32);
                \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.6\ := to_unsigned(0, 16);
                \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.7\ := false;
                \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.8\ := to_unsigned(0, 16);
                \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.9\ := to_unsigned(0, 16);
                \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.10\ := to_unsigned(0, 16);
                \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.11\ := to_unsigned(0, 16);
            else 
                case \BitMask::GetMostSignificantOnePosition().0._State\ is 
                    when \BitMask::GetMostSignificantOnePosition().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\BitMask::GetMostSignificantOnePosition().0._Started\ = true) then 
                            \BitMask::GetMostSignificantOnePosition().0._State\ := \BitMask::GetMostSignificantOnePosition().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::GetMostSignificantOnePosition().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\BitMask::GetMostSignificantOnePosition().0._Started\ = true) then 
                            \BitMask::GetMostSignificantOnePosition().0._Finished\ <= true;
                        else 
                            \BitMask::GetMostSignificantOnePosition().0._Finished\ <= false;
                            \BitMask::GetMostSignificantOnePosition().0._State\ := \BitMask::GetMostSignificantOnePosition().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::GetMostSignificantOnePosition().0._State_2\ => 
                        \BitMask::GetMostSignificantOnePosition().0.this\ := \BitMask::GetMostSignificantOnePosition().0.this.parameter.In\;
                        \BitMask::GetMostSignificantOnePosition().0.num\ := to_unsigned(0, 16);
                        \BitMask::GetMostSignificantOnePosition().0.num2\ := to_unsigned(1, 16);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.0\ := \BitMask::GetMostSignificantOnePosition().0.num2\ <= \BitMask::GetMostSignificantOnePosition().0.this\.\SegmentCount\;
                        if (\BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.0\) then 
                            \BitMask::GetMostSignificantOnePosition().0._State\ := \BitMask::GetMostSignificantOnePosition().0._State_3\;
                        else 
                            \BitMask::GetMostSignificantOnePosition().0._State\ := \BitMask::GetMostSignificantOnePosition().0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::GetMostSignificantOnePosition().0._State_3\ => 
                        -- Repeated state of the while loop which was started in state \BitMask::GetMostSignificantOnePosition().0._State_2\.
                        -- The while loop's condition:
                        \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.1\ := \BitMask::GetMostSignificantOnePosition().0.num2\ <= \BitMask::GetMostSignificantOnePosition().0.this\.\SegmentCount\;
                        if (\BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.1\) then 
                            \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.2\ := resize(signed(\BitMask::GetMostSignificantOnePosition().0.this\.\SegmentCount\ - \BitMask::GetMostSignificantOnePosition().0.num2\), 32);
                            \BitMask::GetMostSignificantOnePosition().0.num3\ := \BitMask::GetMostSignificantOnePosition().0.this\.\Segments\(to_integer((\BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.2\)));
                            -- Starting a while loop.
                            -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                            \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.3\ := \BitMask::GetMostSignificantOnePosition().0.num3\ > to_unsigned(0, 32);
                            if (\BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.3\) then 
                                \BitMask::GetMostSignificantOnePosition().0._State\ := \BitMask::GetMostSignificantOnePosition().0._State_5\;
                            else 
                                \BitMask::GetMostSignificantOnePosition().0._State\ := \BitMask::GetMostSignificantOnePosition().0._State_6\;
                            end if;
                        else 
                            \BitMask::GetMostSignificantOnePosition().0._State\ := \BitMask::GetMostSignificantOnePosition().0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \BitMask::GetMostSignificantOnePosition().0._State_4\ => 
                        -- State after the while loop which was started in state \BitMask::GetMostSignificantOnePosition().0._State_2\.
                        \BitMask::GetMostSignificantOnePosition().0.result\ := to_unsigned(0, 16);
                        \BitMask::GetMostSignificantOnePosition().0.return\ <= to_unsigned(0, 16);
                        \BitMask::GetMostSignificantOnePosition().0._State\ := \BitMask::GetMostSignificantOnePosition().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::GetMostSignificantOnePosition().0._State_5\ => 
                        -- Repeated state of the while loop which was started in state \BitMask::GetMostSignificantOnePosition().0._State_3\.
                        -- The while loop's condition:
                        \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.4\ := \BitMask::GetMostSignificantOnePosition().0.num3\ > to_unsigned(0, 32);
                        if (\BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.4\) then 
                            \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.5\ := shift_right(\BitMask::GetMostSignificantOnePosition().0.num3\, to_integer(to_signed(1, 32)));
                            \BitMask::GetMostSignificantOnePosition().0.num3\ := \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.5\;
                            \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.6\ := \BitMask::GetMostSignificantOnePosition().0.num\ + to_unsigned(1, 16);
                            \BitMask::GetMostSignificantOnePosition().0.num\ := \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.6\;
                            \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.7\ := \BitMask::GetMostSignificantOnePosition().0.num3\ = to_unsigned(0, 32);
                            \BitMask::GetMostSignificantOnePosition().0.flag\ := \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.7\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \BitMask::GetMostSignificantOnePosition().0._State_8\ and ends in state \BitMask::GetMostSignificantOnePosition().0._State_8\.
                            --     * Execution after either branch will continue in the following state: \BitMask::GetMostSignificantOnePosition().0._State_7\.

                            if (\BitMask::GetMostSignificantOnePosition().0.flag\) then 
                                \BitMask::GetMostSignificantOnePosition().0._State\ := \BitMask::GetMostSignificantOnePosition().0._State_8\;
                            else 
                                -- There was no false branch, so going directly to the state after the if-else.
                                \BitMask::GetMostSignificantOnePosition().0._State\ := \BitMask::GetMostSignificantOnePosition().0._State_7\;
                            end if;
                        else 
                            \BitMask::GetMostSignificantOnePosition().0._State\ := \BitMask::GetMostSignificantOnePosition().0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.4
                    when \BitMask::GetMostSignificantOnePosition().0._State_6\ => 
                        -- State after the while loop which was started in state \BitMask::GetMostSignificantOnePosition().0._State_3\.
                        \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.11\ := \BitMask::GetMostSignificantOnePosition().0.num2\ + to_unsigned(1, 16);
                        \BitMask::GetMostSignificantOnePosition().0.num2\ := \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.11\;
                        -- Returning to the repeated state of the while loop which was started in state \BitMask::GetMostSignificantOnePosition().0._State_2\ if the loop wasn't exited with a state change.
                        if (\BitMask::GetMostSignificantOnePosition().0._State\ = \BitMask::GetMostSignificantOnePosition().0._State_6\) then 
                            \BitMask::GetMostSignificantOnePosition().0._State\ := \BitMask::GetMostSignificantOnePosition().0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::GetMostSignificantOnePosition().0._State_7\ => 
                        -- State after the if-else which was started in state \BitMask::GetMostSignificantOnePosition().0._State_5\.
                        -- Returning to the repeated state of the while loop which was started in state \BitMask::GetMostSignificantOnePosition().0._State_3\ if the loop wasn't exited with a state change.
                        if (\BitMask::GetMostSignificantOnePosition().0._State\ = \BitMask::GetMostSignificantOnePosition().0._State_7\) then 
                            \BitMask::GetMostSignificantOnePosition().0._State\ := \BitMask::GetMostSignificantOnePosition().0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::GetMostSignificantOnePosition().0._State_8\ => 
                        -- True branch of the if-else started in state \BitMask::GetMostSignificantOnePosition().0._State_5\.
                        \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.8\ := \BitMask::GetMostSignificantOnePosition().0.this\.\SegmentCount\ - \BitMask::GetMostSignificantOnePosition().0.num2\;
                        \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.9\ := resize(\BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.8\ * to_unsigned(32, 16), 16);
                        \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.10\ := \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.9\ + \BitMask::GetMostSignificantOnePosition().0.num\;
                        \BitMask::GetMostSignificantOnePosition().0.result\ := \BitMask::GetMostSignificantOnePosition().0.binaryOperationResult.10\;
                        \BitMask::GetMostSignificantOnePosition().0.return\ <= \BitMask::GetMostSignificantOnePosition().0.result\;
                        \BitMask::GetMostSignificantOnePosition().0._State\ := \BitMask::GetMostSignificantOnePosition().0._State_1\;
                        -- Going to the state after the if-else which was started in state \BitMask::GetMostSignificantOnePosition().0._State_5\.
                        if (\BitMask::GetMostSignificantOnePosition().0._State\ = \BitMask::GetMostSignificantOnePosition().0._State_8\) then 
                            \BitMask::GetMostSignificantOnePosition().0._State\ := \BitMask::GetMostSignificantOnePosition().0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                end case;
            end if;
        end if;
    end process;
    -- System.UInt16 Lombiq.Unum.BitMask::GetMostSignificantOnePosition().0 state machine end


    -- System.UInt16 Lombiq.Unum.BitMask::GetLeastSignificantOnePosition().0 state machine start
    \BitMask::GetLeastSignificantOnePosition().0._StateMachine\: process (\Clock\) 
        Variable \BitMask::GetLeastSignificantOnePosition().0._State\: \BitMask::GetLeastSignificantOnePosition().0._States\ := \BitMask::GetLeastSignificantOnePosition().0._State_0\;
        Variable \BitMask::GetLeastSignificantOnePosition().0.this\: \Lombiq.Unum.BitMask\;
        Variable \BitMask::GetLeastSignificantOnePosition().0.num\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::GetLeastSignificantOnePosition().0.num2\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::GetLeastSignificantOnePosition().0.num3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::GetLeastSignificantOnePosition().0.flag\: boolean := false;
        Variable \BitMask::GetLeastSignificantOnePosition().0.flag2\: boolean := false;
        Variable \BitMask::GetLeastSignificantOnePosition().0.result\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.0\: boolean := false;
        Variable \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.1\: boolean := false;
        Variable \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.2\: boolean := false;
        Variable \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.3\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.4\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::GetLeastSignificantOnePosition().0.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.5\: boolean := false;
        Variable \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.6\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::GetLeastSignificantOnePosition().0.clockCyclesWaitedForBinaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.7\: boolean := false;
        Variable \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.8\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.9\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.10\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \BitMask::GetLeastSignificantOnePosition().0.clockCyclesWaitedForBinaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.11\: boolean := false;
        Variable \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.12\: unsigned(15 downto 0) := to_unsigned(0, 16);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \BitMask::GetLeastSignificantOnePosition().0._Finished\ <= false;
                \BitMask::GetLeastSignificantOnePosition().0.return\ <= to_unsigned(0, 16);
                \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_0\;
                \BitMask::GetLeastSignificantOnePosition().0.num\ := to_unsigned(0, 16);
                \BitMask::GetLeastSignificantOnePosition().0.num2\ := to_unsigned(0, 16);
                \BitMask::GetLeastSignificantOnePosition().0.num3\ := to_unsigned(0, 32);
                \BitMask::GetLeastSignificantOnePosition().0.flag\ := false;
                \BitMask::GetLeastSignificantOnePosition().0.flag2\ := false;
                \BitMask::GetLeastSignificantOnePosition().0.result\ := to_unsigned(0, 16);
                \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.0\ := false;
                \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.1\ := false;
                \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.2\ := false;
                \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.3\ := to_unsigned(0, 16);
                \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.4\ := to_unsigned(0, 32);
                \BitMask::GetLeastSignificantOnePosition().0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.5\ := false;
                \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.6\ := to_unsigned(0, 32);
                \BitMask::GetLeastSignificantOnePosition().0.clockCyclesWaitedForBinaryOperationResult.1\ := to_signed(0, 32);
                \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.7\ := false;
                \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.8\ := to_unsigned(0, 16);
                \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.9\ := to_unsigned(0, 32);
                \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.10\ := to_unsigned(0, 32);
                \BitMask::GetLeastSignificantOnePosition().0.clockCyclesWaitedForBinaryOperationResult.2\ := to_signed(0, 32);
                \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.11\ := false;
                \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.12\ := to_unsigned(0, 16);
            else 
                case \BitMask::GetLeastSignificantOnePosition().0._State\ is 
                    when \BitMask::GetLeastSignificantOnePosition().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\BitMask::GetLeastSignificantOnePosition().0._Started\ = true) then 
                            \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::GetLeastSignificantOnePosition().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\BitMask::GetLeastSignificantOnePosition().0._Started\ = true) then 
                            \BitMask::GetLeastSignificantOnePosition().0._Finished\ <= true;
                        else 
                            \BitMask::GetLeastSignificantOnePosition().0._Finished\ <= false;
                            \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::GetLeastSignificantOnePosition().0._State_2\ => 
                        \BitMask::GetLeastSignificantOnePosition().0.this\ := \BitMask::GetLeastSignificantOnePosition().0.this.parameter.In\;
                        \BitMask::GetLeastSignificantOnePosition().0.num\ := to_unsigned(1, 16);
                        \BitMask::GetLeastSignificantOnePosition().0.num2\ := to_unsigned(0, 16);
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.0\ := \BitMask::GetLeastSignificantOnePosition().0.num2\ < \BitMask::GetLeastSignificantOnePosition().0.this\.\SegmentCount\;
                        if (\BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.0\) then 
                            \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_3\;
                        else 
                            \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::GetLeastSignificantOnePosition().0._State_3\ => 
                        -- Repeated state of the while loop which was started in state \BitMask::GetLeastSignificantOnePosition().0._State_2\.
                        -- The while loop's condition:
                        \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.1\ := \BitMask::GetLeastSignificantOnePosition().0.num2\ < \BitMask::GetLeastSignificantOnePosition().0.this\.\SegmentCount\;
                        if (\BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.1\) then 
                            \BitMask::GetLeastSignificantOnePosition().0.num3\ := \BitMask::GetLeastSignificantOnePosition().0.this\.\Segments\(to_integer(resize(signed(\BitMask::GetLeastSignificantOnePosition().0.num2\), 32)));
                            \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.2\ := \BitMask::GetLeastSignificantOnePosition().0.num3\ = to_unsigned(0, 32);
                            \BitMask::GetLeastSignificantOnePosition().0.flag\ := \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.2\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \BitMask::GetLeastSignificantOnePosition().0._State_6\ and ends in state \BitMask::GetLeastSignificantOnePosition().0._State_6\.
                            --     * The false branch starts in state \BitMask::GetLeastSignificantOnePosition().0._State_7\ and ends in state \BitMask::GetLeastSignificantOnePosition().0._State_16\.
                            --     * Execution after either branch will continue in the following state: \BitMask::GetLeastSignificantOnePosition().0._State_5\.

                            if (\BitMask::GetLeastSignificantOnePosition().0.flag\) then 
                                \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_6\;
                            else 
                                \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_7\;
                            end if;
                        else 
                            \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \BitMask::GetLeastSignificantOnePosition().0._State_4\ => 
                        -- State after the while loop which was started in state \BitMask::GetLeastSignificantOnePosition().0._State_2\.
                        \BitMask::GetLeastSignificantOnePosition().0.result\ := to_unsigned(0, 16);
                        \BitMask::GetLeastSignificantOnePosition().0.return\ <= to_unsigned(0, 16);
                        \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::GetLeastSignificantOnePosition().0._State_5\ => 
                        -- State after the if-else which was started in state \BitMask::GetLeastSignificantOnePosition().0._State_3\.
                        \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.12\ := \BitMask::GetLeastSignificantOnePosition().0.num2\ + to_unsigned(1, 16);
                        \BitMask::GetLeastSignificantOnePosition().0.num2\ := \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.12\;
                        -- Returning to the repeated state of the while loop which was started in state \BitMask::GetLeastSignificantOnePosition().0._State_2\ if the loop wasn't exited with a state change.
                        if (\BitMask::GetLeastSignificantOnePosition().0._State\ = \BitMask::GetLeastSignificantOnePosition().0._State_5\) then 
                            \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::GetLeastSignificantOnePosition().0._State_6\ => 
                        -- True branch of the if-else started in state \BitMask::GetLeastSignificantOnePosition().0._State_3\.
                        \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.3\ := \BitMask::GetLeastSignificantOnePosition().0.num\ + to_unsigned(32, 16);
                        \BitMask::GetLeastSignificantOnePosition().0.num\ := \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.3\;
                        -- Going to the state after the if-else which was started in state \BitMask::GetLeastSignificantOnePosition().0._State_3\.
                        if (\BitMask::GetLeastSignificantOnePosition().0._State\ = \BitMask::GetLeastSignificantOnePosition().0._State_6\) then 
                            \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::GetLeastSignificantOnePosition().0._State_7\ => 
                        -- False branch of the if-else started in state \BitMask::GetLeastSignificantOnePosition().0._State_3\.
                        -- Starting a while loop.
                        -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                        \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_10\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::GetLeastSignificantOnePosition().0._State_8\ => 
                        -- Repeated state of the while loop which was started in state \BitMask::GetLeastSignificantOnePosition().0._State_7\.
                        -- The while loop's condition:
                        \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_12\;
                        if (\BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.7\) then 
                            \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.8\ := \BitMask::GetLeastSignificantOnePosition().0.num\ + to_unsigned(1, 16);
                            \BitMask::GetLeastSignificantOnePosition().0.num\ := \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.8\;
                            \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.9\ := shift_right(\BitMask::GetLeastSignificantOnePosition().0.num3\, to_integer(to_signed(1, 32)));
                            \BitMask::GetLeastSignificantOnePosition().0.num3\ := \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.9\;
                            -- Returning to the repeated state of the while loop which was started in state \BitMask::GetLeastSignificantOnePosition().0._State_7\ if the loop wasn't exited with a state change.
                            if (\BitMask::GetLeastSignificantOnePosition().0._State\ = \BitMask::GetLeastSignificantOnePosition().0._State_13\) then 
                                \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_8\;
                            end if;
                        else 
                            \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_9\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::GetLeastSignificantOnePosition().0._State_9\ => 
                        -- State after the while loop which was started in state \BitMask::GetLeastSignificantOnePosition().0._State_7\.
                        \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_14\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::GetLeastSignificantOnePosition().0._State_10\ => 
                        -- Waiting for the result to appear in \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.4\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\BitMask::GetLeastSignificantOnePosition().0.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_11\;
                            \BitMask::GetLeastSignificantOnePosition().0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \BitMask::GetLeastSignificantOnePosition().0.clockCyclesWaitedForBinaryOperationResult.0\ := \BitMask::GetLeastSignificantOnePosition().0.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.4\ := \BitMask::GetLeastSignificantOnePosition().0.num3\ mod to_unsigned(2, 32);
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \BitMask::GetLeastSignificantOnePosition().0._State_11\ => 
                        \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.5\ := \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.4\ = to_unsigned(0, 32);
                        if (\BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.5\) then 
                            \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_8\;
                        else 
                            \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_9\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::GetLeastSignificantOnePosition().0._State_12\ => 
                        -- Waiting for the result to appear in \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.6\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\BitMask::GetLeastSignificantOnePosition().0.clockCyclesWaitedForBinaryOperationResult.1\ >= to_signed(7, 32)) then 
                            \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_13\;
                            \BitMask::GetLeastSignificantOnePosition().0.clockCyclesWaitedForBinaryOperationResult.1\ := to_signed(0, 32);
                        else 
                            \BitMask::GetLeastSignificantOnePosition().0.clockCyclesWaitedForBinaryOperationResult.1\ := \BitMask::GetLeastSignificantOnePosition().0.clockCyclesWaitedForBinaryOperationResult.1\ + to_signed(1, 32);
                        end if;
                        \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.6\ := \BitMask::GetLeastSignificantOnePosition().0.num3\ mod to_unsigned(2, 32);
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \BitMask::GetLeastSignificantOnePosition().0._State_13\ => 
                        \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.7\ := \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.6\ = to_unsigned(0, 32);
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \BitMask::GetLeastSignificantOnePosition().0._State_14\ => 
                        -- Waiting for the result to appear in \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.10\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\BitMask::GetLeastSignificantOnePosition().0.clockCyclesWaitedForBinaryOperationResult.2\ >= to_signed(7, 32)) then 
                            \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_15\;
                            \BitMask::GetLeastSignificantOnePosition().0.clockCyclesWaitedForBinaryOperationResult.2\ := to_signed(0, 32);
                        else 
                            \BitMask::GetLeastSignificantOnePosition().0.clockCyclesWaitedForBinaryOperationResult.2\ := \BitMask::GetLeastSignificantOnePosition().0.clockCyclesWaitedForBinaryOperationResult.2\ + to_signed(1, 32);
                        end if;
                        \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.10\ := \BitMask::GetLeastSignificantOnePosition().0.num3\ mod to_unsigned(2, 32);
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \BitMask::GetLeastSignificantOnePosition().0._State_15\ => 
                        \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.11\ := \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.10\ = to_unsigned(1, 32);
                        \BitMask::GetLeastSignificantOnePosition().0.flag2\ := \BitMask::GetLeastSignificantOnePosition().0.binaryOperationResult.11\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \BitMask::GetLeastSignificantOnePosition().0._State_17\ and ends in state \BitMask::GetLeastSignificantOnePosition().0._State_17\.
                        --     * Execution after either branch will continue in the following state: \BitMask::GetLeastSignificantOnePosition().0._State_16\.

                        if (\BitMask::GetLeastSignificantOnePosition().0.flag2\) then 
                            \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_17\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_16\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \BitMask::GetLeastSignificantOnePosition().0._State_16\ => 
                        -- State after the if-else which was started in state \BitMask::GetLeastSignificantOnePosition().0._State_15\.
                        -- Going to the state after the if-else which was started in state \BitMask::GetLeastSignificantOnePosition().0._State_3\.
                        if (\BitMask::GetLeastSignificantOnePosition().0._State\ = \BitMask::GetLeastSignificantOnePosition().0._State_16\) then 
                            \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::GetLeastSignificantOnePosition().0._State_17\ => 
                        -- True branch of the if-else started in state \BitMask::GetLeastSignificantOnePosition().0._State_15\.
                        \BitMask::GetLeastSignificantOnePosition().0.result\ := \BitMask::GetLeastSignificantOnePosition().0.num\;
                        \BitMask::GetLeastSignificantOnePosition().0.return\ <= \BitMask::GetLeastSignificantOnePosition().0.result\;
                        \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_1\;
                        -- Going to the state after the if-else which was started in state \BitMask::GetLeastSignificantOnePosition().0._State_15\.
                        if (\BitMask::GetLeastSignificantOnePosition().0._State\ = \BitMask::GetLeastSignificantOnePosition().0._State_17\) then 
                            \BitMask::GetLeastSignificantOnePosition().0._State\ := \BitMask::GetLeastSignificantOnePosition().0._State_16\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.UInt16 Lombiq.Unum.BitMask::GetLeastSignificantOnePosition().0 state machine end


    -- System.UInt32 Lombiq.Unum.BitMask::GetLowest32Bits().0 state machine start
    \BitMask::GetLowest32Bits().0._StateMachine\: process (\Clock\) 
        Variable \BitMask::GetLowest32Bits().0._State\: \BitMask::GetLowest32Bits().0._States\ := \BitMask::GetLowest32Bits().0._State_0\;
        Variable \BitMask::GetLowest32Bits().0.this\: \Lombiq.Unum.BitMask\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \BitMask::GetLowest32Bits().0._Finished\ <= false;
                \BitMask::GetLowest32Bits().0.return\ <= to_unsigned(0, 32);
                \BitMask::GetLowest32Bits().0._State\ := \BitMask::GetLowest32Bits().0._State_0\;
            else 
                case \BitMask::GetLowest32Bits().0._State\ is 
                    when \BitMask::GetLowest32Bits().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\BitMask::GetLowest32Bits().0._Started\ = true) then 
                            \BitMask::GetLowest32Bits().0._State\ := \BitMask::GetLowest32Bits().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::GetLowest32Bits().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\BitMask::GetLowest32Bits().0._Started\ = true) then 
                            \BitMask::GetLowest32Bits().0._Finished\ <= true;
                        else 
                            \BitMask::GetLowest32Bits().0._Finished\ <= false;
                            \BitMask::GetLowest32Bits().0._State\ := \BitMask::GetLowest32Bits().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \BitMask::GetLowest32Bits().0._State_2\ => 
                        \BitMask::GetLowest32Bits().0.this\ := \BitMask::GetLowest32Bits().0.this.parameter.In\;
                        \BitMask::GetLowest32Bits().0.return\ <= \BitMask::GetLowest32Bits().0.this\.\Segments\(to_integer(to_signed(0, 32)));
                        \BitMask::GetLowest32Bits().0._State\ := \BitMask::GetLowest32Bits().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.UInt32 Lombiq.Unum.BitMask::GetLowest32Bits().0 state machine end


    -- System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment).0 state machine start
    \Unum::.ctor(UnumEnvironment).0._StateMachine\: process (\Clock\) 
        Variable \Unum::.ctor(UnumEnvironment).0._State\: \Unum::.ctor(UnumEnvironment).0._States\ := \Unum::.ctor(UnumEnvironment).0._State_0\;
        Variable \Unum::.ctor(UnumEnvironment).0.this\: \Lombiq.Unum.Unum\;
        Variable \Unum::.ctor(UnumEnvironment).0.environment\: \Lombiq.Unum.UnumEnvironment\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::.ctor(UnumEnvironment).0._Finished\ <= false;
                \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\ <= false;
                \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= false;
                \Unum::.ctor(UnumEnvironment).0._State\ := \Unum::.ctor(UnumEnvironment).0._State_0\;
            else 
                case \Unum::.ctor(UnumEnvironment).0._State\ is 
                    when \Unum::.ctor(UnumEnvironment).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::.ctor(UnumEnvironment).0._Started\ = true) then 
                            \Unum::.ctor(UnumEnvironment).0._State\ := \Unum::.ctor(UnumEnvironment).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::.ctor(UnumEnvironment).0._Started\ = true) then 
                            \Unum::.ctor(UnumEnvironment).0._Finished\ <= true;
                        else 
                            \Unum::.ctor(UnumEnvironment).0._Finished\ <= false;
                            \Unum::.ctor(UnumEnvironment).0._State\ := \Unum::.ctor(UnumEnvironment).0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \Unum::.ctor(UnumEnvironment).0.this.parameter.Out\ <= \Unum::.ctor(UnumEnvironment).0.this\;
                        \Unum::.ctor(UnumEnvironment).0.environment.parameter.Out\ <= \Unum::.ctor(UnumEnvironment).0.environment\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment).0._State_2\ => 
                        \Unum::.ctor(UnumEnvironment).0.this\ := \Unum::.ctor(UnumEnvironment).0.this.parameter.In\;
                        \Unum::.ctor(UnumEnvironment).0.environment\ := \Unum::.ctor(UnumEnvironment).0.environment.parameter.In\;
                        \Unum::.ctor(UnumEnvironment).0.this\.\_environment\ := \Unum::.ctor(UnumEnvironment).0.environment\;
                        -- Initializing record fields to their defaults.
                        \Unum::.ctor(UnumEnvironment).0.this\.\UnumBits\.\IsNull\ := false;
                        \Unum::.ctor(UnumEnvironment).0.this\.\UnumBits\.\Size\ := to_unsigned(0, 16);
                        \Unum::.ctor(UnumEnvironment).0.this\.\UnumBits\.\SegmentCount\ := to_unsigned(0, 16);
                        \Unum::.ctor(UnumEnvironment).0.this\.\UnumBits\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                        \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment).0.this\.\UnumBits\;
                        \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment).0.this\.\_environment\.\Size\;
                        \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\ <= False;
                        \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= true;
                        \Unum::.ctor(UnumEnvironment).0._State\ := \Unum::.ctor(UnumEnvironment).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment).0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                        if (\Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ = \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\) then 
                            \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= false;
                            \Unum::.ctor(UnumEnvironment).0.this\.\UnumBits\ := \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\;
                            \Unum::.ctor(UnumEnvironment).0._State\ := \Unum::.ctor(UnumEnvironment).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment).0 state machine end


    -- System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,Lombiq.Unum.BitMask).0 state machine start
    \Unum::.ctor(UnumEnvironment,BitMask).0._StateMachine\: process (\Clock\) 
        Variable \Unum::.ctor(UnumEnvironment,BitMask).0._State\: \Unum::.ctor(UnumEnvironment,BitMask).0._States\ := \Unum::.ctor(UnumEnvironment,BitMask).0._State_0\;
        Variable \Unum::.ctor(UnumEnvironment,BitMask).0.this\: \Lombiq.Unum.Unum\;
        Variable \Unum::.ctor(UnumEnvironment,BitMask).0.environment\: \Lombiq.Unum.UnumEnvironment\;
        Variable \Unum::.ctor(UnumEnvironment,BitMask).0.bits\: \Lombiq.Unum.BitMask\;
        Variable \Unum::.ctor(UnumEnvironment,BitMask).0.return.0\: \Lombiq.Unum.BitMask\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::.ctor(UnumEnvironment,BitMask).0._Finished\ <= false;
                \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 32));
                \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Started.0\ <= false;
                \Unum::.ctor(UnumEnvironment,BitMask).0._State\ := \Unum::.ctor(UnumEnvironment,BitMask).0._State_0\;
            else 
                case \Unum::.ctor(UnumEnvironment,BitMask).0._State\ is 
                    when \Unum::.ctor(UnumEnvironment,BitMask).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::.ctor(UnumEnvironment,BitMask).0._Started\ = true) then 
                            \Unum::.ctor(UnumEnvironment,BitMask).0._State\ := \Unum::.ctor(UnumEnvironment,BitMask).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,BitMask).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::.ctor(UnumEnvironment,BitMask).0._Started\ = true) then 
                            \Unum::.ctor(UnumEnvironment,BitMask).0._Finished\ <= true;
                        else 
                            \Unum::.ctor(UnumEnvironment,BitMask).0._Finished\ <= false;
                            \Unum::.ctor(UnumEnvironment,BitMask).0._State\ := \Unum::.ctor(UnumEnvironment,BitMask).0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \Unum::.ctor(UnumEnvironment,BitMask).0.this.parameter.Out\ <= \Unum::.ctor(UnumEnvironment,BitMask).0.this\;
                        \Unum::.ctor(UnumEnvironment,BitMask).0.environment.parameter.Out\ <= \Unum::.ctor(UnumEnvironment,BitMask).0.environment\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,BitMask).0._State_2\ => 
                        \Unum::.ctor(UnumEnvironment,BitMask).0.this\ := \Unum::.ctor(UnumEnvironment,BitMask).0.this.parameter.In\;
                        \Unum::.ctor(UnumEnvironment,BitMask).0.environment\ := \Unum::.ctor(UnumEnvironment,BitMask).0.environment.parameter.In\;
                        \Unum::.ctor(UnumEnvironment,BitMask).0.bits\ := \Unum::.ctor(UnumEnvironment,BitMask).0.bits.parameter.In\;
                        \Unum::.ctor(UnumEnvironment,BitMask).0.this\.\_environment\ := \Unum::.ctor(UnumEnvironment,BitMask).0.environment\;
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::FromImmutableArray(System.UInt32[],System.UInt16)
                        \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16).segments.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,BitMask).0.bits\.\Segments\;
                        \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16).size.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,BitMask).0.this\.\_environment\.\Size\;
                        \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Started.0\ <= true;
                        \Unum::.ctor(UnumEnvironment,BitMask).0._State\ := \Unum::.ctor(UnumEnvironment,BitMask).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,BitMask).0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::FromImmutableArray(System.UInt32[],System.UInt16)
                        if (\Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Started.0\ = \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Finished.0\) then 
                            \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Started.0\ <= false;
                            \Unum::.ctor(UnumEnvironment,BitMask).0.return.0\ := \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16).return.0\;
                            \Unum::.ctor(UnumEnvironment,BitMask).0.bits\.\Segments\ := \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16).segments.parameter.In.0\;
                            \Unum::.ctor(UnumEnvironment,BitMask).0.this\.\UnumBits\ := \Unum::.ctor(UnumEnvironment,BitMask).0.return.0\;
                            \Unum::.ctor(UnumEnvironment,BitMask).0._State\ := \Unum::.ctor(UnumEnvironment,BitMask).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,Lombiq.Unum.BitMask).0 state machine end


    -- System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.UInt32[],System.Boolean).0 state machine start
    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._StateMachine\: process (\Clock\) 
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\: \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._States\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_0\;
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.this\: \Lombiq.Unum.Unum\;
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.environment\: \Lombiq.Unum.UnumEnvironment\;
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.value\: \unsigned32_Array\(0 to 0) := (others => to_unsigned(0, 32));
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.negative\: boolean := false;
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.flag\: boolean := false;
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.exponent\: \Lombiq.Unum.BitMask\;
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.left\: \Lombiq.Unum.BitMask\;
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.num\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.flag2\: boolean := false;
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.right\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.fraction\: \Lombiq.Unum.BitMask\;
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.num2\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.flag3\: boolean := false;
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.0\: boolean := false;
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.1\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.arraye795bd01e461b0dce534a453220c7f445988b9bd9f9fb443b451fcbaf1ac12a0\: \unsigned32_Array\(0 to 0) := (others => to_unsigned(0, 32));
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.2\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.3\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.4\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.5\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.6\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.3\: boolean := false;
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.4\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.5\: boolean := false;
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.6\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.7\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.8\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.7\: \Lombiq.Unum.BitMask\;
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.8\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.9\: \Lombiq.Unum.BitMask\;
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.10\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.11\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.9\: boolean := false;
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.10\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.12\: \Lombiq.Unum.BitMask\;
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.conditional1059d8789965c7346ddefe992fa75edc6265395c1804dfe1295a035696e9157b\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.11\: boolean := false;
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.12\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.conditional11166ff980773138629b8148bc5ab3129946c943a4d67b94f55ae0052361c700\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.13\: boolean := false;
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.14\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.13\: \Lombiq.Unum.BitMask\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._Finished\ <= false;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.value.parameter.Out\ <= (others => to_unsigned(0, 32));
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 32));
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ <= false;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size()._Started.0\ <= false;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition()._Started.0\ <= false;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits()._Started.0\ <= false;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\ <= to_unsigned(0, 32);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ <= false;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::ShiftOutLeastSignificantZeros()._Started.0\ <= false;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::SetZero(UInt16).index.parameter.Out.0\ <= to_unsigned(0, 16);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::SetZero(UInt16)._Started.0\ <= false;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).signBit.parameter.Out.0\ <= false;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).uncertainityBit.parameter.Out.0\ <= false;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).exponentSize.parameter.Out.0\ <= to_unsigned(0, 8);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).fractionSize.parameter.Out.0\ <= to_unsigned(0, 16);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Started.0\ <= false;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_0\;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.value\ := (others => to_unsigned(0, 32));
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.negative\ := false;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.flag\ := false;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.num\ := to_unsigned(0, 16);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.flag2\ := false;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.right\ := to_signed(0, 32);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.num2\ := to_unsigned(0, 16);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.flag3\ := false;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.0\ := false;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.1\ := to_unsigned(0, 16);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.arraye795bd01e461b0dce534a453220c7f445988b9bd9f9fb443b451fcbaf1ac12a0\ := (others => to_unsigned(0, 32));
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.2\ := to_unsigned(0, 16);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.0\ := to_unsigned(0, 32);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.3\ := to_unsigned(0, 16);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.4\ := to_unsigned(0, 16);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.5\ := to_unsigned(0, 32);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.6\ := to_unsigned(0, 32);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.1\ := to_unsigned(0, 32);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.2\ := to_unsigned(0, 32);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.3\ := false;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.4\ := to_unsigned(0, 16);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.5\ := false;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.6\ := to_signed(0, 32);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.7\ := to_signed(0, 32);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.8\ := to_signed(0, 32);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.8\ := to_unsigned(0, 16);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.10\ := to_unsigned(0, 16);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.11\ := to_unsigned(0, 32);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.9\ := false;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.10\ := to_unsigned(0, 16);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.conditional1059d8789965c7346ddefe992fa75edc6265395c1804dfe1295a035696e9157b\ := to_unsigned(0, 16);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.11\ := false;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.12\ := to_unsigned(0, 16);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.conditional11166ff980773138629b8148bc5ab3129946c943a4d67b94f55ae0052361c700\ := to_unsigned(0, 16);
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.13\ := false;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.14\ := to_unsigned(0, 16);
            else 
                case \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ is 
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._Started\ = true) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._Started\ = true) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._Finished\ <= true;
                        else 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._Finished\ <= false;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.this.parameter.Out\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.this\;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.environment.parameter.Out\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.environment\;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.value.parameter.Out\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.value\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_2\ => 
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.this\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.this.parameter.In\;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.environment\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.environment.parameter.In\;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.value\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.value.parameter.In\;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.negative\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.negative.parameter.In\;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.this\.\_environment\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.environment\;
                        -- Initializing record fields to their defaults.
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.this\.\UnumBits\.\IsNull\ := false;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.this\.\UnumBits\.\Size\ := to_unsigned(0, 16);
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.this\.\UnumBits\.\SegmentCount\ := to_unsigned(0, 16);
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.this\.\UnumBits\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.this\.\UnumBits\;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\(0 to 0) <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.value\;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.environment\.\Size\;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= true;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.this\.\UnumBits\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.value\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\(0 to 0);
                            -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.BitMask::op_Equality(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Equality(BitMask,BitMask).left.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.this\.\UnumBits\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Equality(BitMask,BitMask).right.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.this\.\_environment\.\EmptyBitMask\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ <= true;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.BitMask::op_Equality(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ <= false;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.0\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Equality(BitMask,BitMask).return.0\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.flag\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.0\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_6\ and ends in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_37\.
                            --     * Execution after either branch will continue in the following state: \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_5\.

                            if (not(\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.flag\)) then 
                                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_6\;
                            else 
                                -- There was no false branch, so going directly to the state after the if-else.
                                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_5\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_5\ => 
                        -- State after the if-else which was started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_4\.
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_6\ => 
                        -- True branch of the if-else started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_4\.
                        -- Initializing record fields to their defaults.
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.exponent\.\IsNull\ := false;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.exponent\.\Size\ := to_unsigned(0, 16);
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.exponent\.\SegmentCount\ := to_unsigned(0, 16);
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.exponent\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::get_Size()
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size().this.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.this\;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size()._Started.0\ <= true;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_7\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_7\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::get_Size()
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size()._Started.0\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size()._Finished.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size()._Started.0\ <= false;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.1\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size().return.0\;
                            -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.exponent\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\(0 to 0) <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.value\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.1\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= true;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_8\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.exponent\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.value\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\(0 to 0);
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.arraye795bd01e461b0dce534a453220c7f445988b9bd9f9fb443b451fcbaf1ac12a0\ := (others => to_unsigned(0, 32));
                            -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.BitMask::GetMostSignificantOnePosition()
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition().this.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.exponent\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition()._Started.0\ <= true;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_9\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_9\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.BitMask::GetMostSignificantOnePosition()
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition()._Started.0\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition()._Finished.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition()._Started.0\ <= false;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.2\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition().return.0\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.0\ := resize(\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.2\ - to_unsigned(1, 16), 32);
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.arraye795bd01e461b0dce534a453220c7f445988b9bd9f9fb443b451fcbaf1ac12a0\(to_integer(to_signed(0, 32))) := (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.0\);
                            -- Initializing record fields to their defaults.
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.left\.\IsNull\ := false;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.left\.\Size\ := to_unsigned(0, 16);
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.left\.\SegmentCount\ := to_unsigned(0, 16);
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.left\.\Segments\ := (others => to_unsigned(0, 32));
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::get_Size()
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size().this.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.this\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size()._Started.0\ <= true;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_10\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_10\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::get_Size()
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size()._Started.0\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size()._Finished.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size()._Started.0\ <= false;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.3\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size().return.0\;
                            -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.left\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\(0 to 0) <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.arraye795bd01e461b0dce534a453220c7f445988b9bd9f9fb443b451fcbaf1ac12a0\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.3\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= true;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_11\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_11\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.left\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.arraye795bd01e461b0dce534a453220c7f445988b9bd9f9fb443b451fcbaf1ac12a0\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\(0 to 0);
                            -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.BitMask::GetMostSignificantOnePosition()
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition().this.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.left\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition()._Started.0\ <= true;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_12\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_12\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.BitMask::GetMostSignificantOnePosition()
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition()._Started.0\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition()._Finished.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition()._Started.0\ <= false;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.4\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition().return.0\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.num\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.4\;
                            -- Starting state machine invocation for the following method: System.UInt32 Lombiq.Unum.BitMask::GetLowest32Bits()
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits().this.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.left\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits()._Started.0\ <= true;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_13\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_13\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Lombiq.Unum.BitMask::GetLowest32Bits()
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits()._Started.0\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits()._Finished.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits()._Started.0\ <= false;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.5\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits().return.0\;
                            -- The last invocation for the target state machine just finished, so need to start the next one in a later state.
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_14\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_14\ => 
                        -- This state was just added to leave time for the invocation proxy to register that the previous invocation finished.
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_15\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_15\ => 
                        -- Starting state machine invocation for the following method: System.UInt32 Lombiq.Unum.BitMask::GetLowest32Bits()
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits().this.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.left\;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits()._Started.0\ <= true;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_16\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_16\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Lombiq.Unum.BitMask::GetLowest32Bits()
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits()._Started.0\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits()._Finished.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits()._Started.0\ <= false;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.6\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits().return.0\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.1\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.6\ - to_unsigned(1, 32);
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.2\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.5\ and \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.1\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.3\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.2\ > to_unsigned(0, 32);
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.flag2\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.3\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_18\ and ends in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_18\.
                            --     * Execution after either branch will continue in the following state: \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_17\.

                            if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.flag2\) then 
                                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_18\;
                            else 
                                -- There was no false branch, so going directly to the state after the if-else.
                                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_17\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_17\ => 
                        -- State after the if-else which was started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_16\.
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.5\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.num\ = to_unsigned(0, 16);

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_20\ and ends in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_20\.
                        --     * The false branch starts in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_21\ and ends in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_21\.
                        --     * Execution after either branch will continue in the following state: \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_19\.

                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.5\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_20\;
                        else 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_21\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_18\ => 
                        -- True branch of the if-else started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_16\.
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.4\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.num\ + to_unsigned(1, 16);
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.num\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.4\;
                        -- Going to the state after the if-else which was started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_16\.
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_18\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_17\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_19\ => 
                        -- State after the if-else which was started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_17\.
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,System.UInt32)
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Addition(BitMask,UInt32).left.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.left\;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\ <= unsigned(\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.right\);
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ <= true;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_22\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_20\ => 
                        -- True branch of the if-else started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_17\.
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.right\ := to_signed(0, 32);
                        -- Going to the state after the if-else which was started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_17\.
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_20\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_19\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_21\ => 
                        -- False branch of the if-else started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_17\.
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.6\ := resize(signed(\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.num\ - to_unsigned(1, 16)), 32);
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.7\ := resize(shift_left(to_signed(1, 32), to_integer((\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.6\))), 32);
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.8\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.7\ - to_signed(1, 32);
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.right\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.8\;
                        -- Going to the state after the if-else which was started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_17\.
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_21\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_19\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_22\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,System.UInt32)
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ <= false;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.7\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Addition(BitMask,UInt32).return.0\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.exponent\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.7\;
                            -- Initializing record fields to their defaults.
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.fraction\.\IsNull\ := false;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.fraction\.\Size\ := to_unsigned(0, 16);
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.fraction\.\SegmentCount\ := to_unsigned(0, 16);
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.fraction\.\Segments\ := (others => to_unsigned(0, 32));
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::get_Size()
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size().this.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.this\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size()._Started.0\ <= true;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_23\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_23\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::get_Size()
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size()._Started.0\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size()._Finished.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size()._Started.0\ <= false;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.8\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size().return.0\;
                            -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.fraction\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\(0 to 0) <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.value\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.8\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= true;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_24\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_24\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.fraction\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.value\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\(0 to 0);
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::ShiftOutLeastSignificantZeros()
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::ShiftOutLeastSignificantZeros().this.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.fraction\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::ShiftOutLeastSignificantZeros()._Started.0\ <= true;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_25\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_25\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::ShiftOutLeastSignificantZeros()
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::ShiftOutLeastSignificantZeros()._Started.0\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::ShiftOutLeastSignificantZeros()._Finished.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::ShiftOutLeastSignificantZeros()._Started.0\ <= false;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.9\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::ShiftOutLeastSignificantZeros().return.0\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.fraction\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.9\;
                            -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.BitMask::GetMostSignificantOnePosition()
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition().this.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.fraction\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition()._Started.0\ <= true;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_26\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_26\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.BitMask::GetMostSignificantOnePosition()
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition()._Started.0\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition()._Finished.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition()._Started.0\ <= false;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.10\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition().return.0\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.num2\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.10\;
                            -- Starting state machine invocation for the following method: System.UInt32 Lombiq.Unum.BitMask::GetLowest32Bits()
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits().this.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.exponent\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits()._Started.0\ <= true;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_27\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_27\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Lombiq.Unum.BitMask::GetLowest32Bits()
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits()._Started.0\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits()._Finished.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits()._Started.0\ <= false;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.11\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits().return.0\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.9\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.11\ > to_unsigned(0, 32);
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.flag3\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.9\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_29\ and ends in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_30\.
                            --     * Execution after either branch will continue in the following state: \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_28\.

                            if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.flag3\) then 
                                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_29\;
                            else 
                                -- There was no false branch, so going directly to the state after the if-else.
                                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_28\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_28\ => 
                        -- State after the if-else which was started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_27\.
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.11\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.num\ > to_unsigned(0, 16);

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_32\ and ends in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_32\.
                        --     * The false branch starts in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_33\ and ends in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_33\.
                        --     * Execution after either branch will continue in the following state: \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_31\.

                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.11\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_32\;
                        else 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_33\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_29\ => 
                        -- True branch of the if-else started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_27\.
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.10\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.num2\ - to_unsigned(1, 16);
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.num2\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.10\;
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetZero(System.UInt16)
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::SetZero(UInt16).this.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.fraction\;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::SetZero(UInt16).index.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.num2\;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::SetZero(UInt16)._Started.0\ <= true;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_30\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_30\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetZero(System.UInt16)
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::SetZero(UInt16)._Started.0\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::SetZero(UInt16)._Finished.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::SetZero(UInt16)._Started.0\ <= false;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.12\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::SetZero(UInt16).return.0\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.fraction\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.12\;
                            -- Going to the state after the if-else which was started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_27\.
                            if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_30\) then 
                                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_28\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_31\ => 
                        -- State after the if-else which was started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_28\.
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.13\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.num2\ > to_unsigned(0, 16);

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_35\ and ends in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_35\.
                        --     * The false branch starts in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_36\ and ends in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_36\.
                        --     * Execution after either branch will continue in the following state: \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_34\.

                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.13\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_35\;
                        else 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_36\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_32\ => 
                        -- True branch of the if-else started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_28\.
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.12\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.num\ - to_unsigned(1, 16);
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.conditional1059d8789965c7346ddefe992fa75edc6265395c1804dfe1295a035696e9157b\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.12\;
                        -- Going to the state after the if-else which was started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_28\.
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_32\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_31\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_33\ => 
                        -- False branch of the if-else started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_28\.
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.conditional1059d8789965c7346ddefe992fa75edc6265395c1804dfe1295a035696e9157b\ := to_unsigned(0, 16);
                        -- Going to the state after the if-else which was started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_28\.
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_33\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_31\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_34\ => 
                        -- State after the if-else which was started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_31\.
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::SetUnumBits(System.Boolean,Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean,System.Byte,System.UInt16)
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).this.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.this\;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).signBit.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.negative\;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).exponent.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.exponent\;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).fraction.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.fraction\;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).uncertainityBit.parameter.Out.0\ <= False;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).exponentSize.parameter.Out.0\ <= resize((\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.conditional1059d8789965c7346ddefe992fa75edc6265395c1804dfe1295a035696e9157b\), 8);
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).fractionSize.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.conditional11166ff980773138629b8148bc5ab3129946c943a4d67b94f55ae0052361c700\;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Started.0\ <= true;
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_37\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_35\ => 
                        -- True branch of the if-else started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_31\.
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.14\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.num2\ - to_unsigned(1, 16);
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.conditional11166ff980773138629b8148bc5ab3129946c943a4d67b94f55ae0052361c700\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.binaryOperationResult.14\;
                        -- Going to the state after the if-else which was started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_31\.
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_35\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_34\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_36\ => 
                        -- False branch of the if-else started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_31\.
                        \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.conditional11166ff980773138629b8148bc5ab3129946c943a4d67b94f55ae0052361c700\ := to_unsigned(0, 16);
                        -- Going to the state after the if-else which was started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_31\.
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_36\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_34\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_37\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::SetUnumBits(System.Boolean,Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean,System.Byte,System.UInt16)
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Started.0\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Finished.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Started.0\ <= false;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.13\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).return.0\;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.this\.\UnumBits\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.return.13\;
                            -- Going to the state after the if-else which was started in state \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_4\.
                            if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ = \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_37\) then 
                                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State\ := \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._State_5\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.UInt32[],System.Boolean).0 state machine end


    -- System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.Int32).0 state machine start
    \Unum::.ctor(UnumEnvironment,Int32).0._StateMachine\: process (\Clock\) 
        Variable \Unum::.ctor(UnumEnvironment,Int32).0._State\: \Unum::.ctor(UnumEnvironment,Int32).0._States\ := \Unum::.ctor(UnumEnvironment,Int32).0._State_0\;
        Variable \Unum::.ctor(UnumEnvironment,Int32).0.this\: \Lombiq.Unum.Unum\;
        Variable \Unum::.ctor(UnumEnvironment,Int32).0.environment\: \Lombiq.Unum.UnumEnvironment\;
        Variable \Unum::.ctor(UnumEnvironment,Int32).0.value\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::.ctor(UnumEnvironment,Int32).0.array33fbc39d577dad5ed6f3add64bb11d85840cbcf74dc3de0631f99002274571ae\: \unsigned32_Array\(0 to 0) := (others => to_unsigned(0, 32));
        Variable \Unum::.ctor(UnumEnvironment,Int32).0.arrayc56f74e3798679843c34bc7afcaef2219b75aeedea3562d19b496a830cfa8fe8\: \unsigned32_Array\(0 to 0) := (others => to_unsigned(0, 32));
        Variable \Unum::.ctor(UnumEnvironment,Int32).0.conditional65ed64d003b02a249ce90498ecf1a8ab72b84c723e77e357f582c5a48bb18fc1\: \Lombiq.Unum.BitMask\;
        Variable \Unum::.ctor(UnumEnvironment,Int32).0.binaryOperationResult.0\: boolean := false;
        Variable \Unum::.ctor(UnumEnvironment,Int32).0.object739e7c0ee2e2d7e2885cba3d8567c7f7fc002803beba2f5f98ae4af41e10ce82\: \Lombiq.Unum.Unum\;
        Variable \Unum::.ctor(UnumEnvironment,Int32).0.object308d6421e1cd9a8ca8e86fd94126f7dddd720821b3965d0d437be91e799be3b9\: \Lombiq.Unum.Unum\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::.ctor(UnumEnvironment,Int32).0._Finished\ <= false;
                \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).value.parameter.Out.0\ <= (others => to_unsigned(0, 32));
                \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).negative.parameter.Out.0\ <= false;
                \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean)._Started.0\ <= false;
                \Unum::.ctor(UnumEnvironment,Int32).0._State\ := \Unum::.ctor(UnumEnvironment,Int32).0._State_0\;
                \Unum::.ctor(UnumEnvironment,Int32).0.value\ := to_signed(0, 32);
                \Unum::.ctor(UnumEnvironment,Int32).0.array33fbc39d577dad5ed6f3add64bb11d85840cbcf74dc3de0631f99002274571ae\ := (others => to_unsigned(0, 32));
                \Unum::.ctor(UnumEnvironment,Int32).0.arrayc56f74e3798679843c34bc7afcaef2219b75aeedea3562d19b496a830cfa8fe8\ := (others => to_unsigned(0, 32));
                \Unum::.ctor(UnumEnvironment,Int32).0.binaryOperationResult.0\ := false;
            else 
                case \Unum::.ctor(UnumEnvironment,Int32).0._State\ is 
                    when \Unum::.ctor(UnumEnvironment,Int32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::.ctor(UnumEnvironment,Int32).0._Started\ = true) then 
                            \Unum::.ctor(UnumEnvironment,Int32).0._State\ := \Unum::.ctor(UnumEnvironment,Int32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,Int32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::.ctor(UnumEnvironment,Int32).0._Started\ = true) then 
                            \Unum::.ctor(UnumEnvironment,Int32).0._Finished\ <= true;
                        else 
                            \Unum::.ctor(UnumEnvironment,Int32).0._Finished\ <= false;
                            \Unum::.ctor(UnumEnvironment,Int32).0._State\ := \Unum::.ctor(UnumEnvironment,Int32).0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \Unum::.ctor(UnumEnvironment,Int32).0.this.parameter.Out\ <= \Unum::.ctor(UnumEnvironment,Int32).0.this\;
                        \Unum::.ctor(UnumEnvironment,Int32).0.environment.parameter.Out\ <= \Unum::.ctor(UnumEnvironment,Int32).0.environment\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,Int32).0._State_2\ => 
                        \Unum::.ctor(UnumEnvironment,Int32).0.this\ := \Unum::.ctor(UnumEnvironment,Int32).0.this.parameter.In\;
                        \Unum::.ctor(UnumEnvironment,Int32).0.environment\ := \Unum::.ctor(UnumEnvironment,Int32).0.environment.parameter.In\;
                        \Unum::.ctor(UnumEnvironment,Int32).0.value\ := \Unum::.ctor(UnumEnvironment,Int32).0.value.parameter.In\;
                        \Unum::.ctor(UnumEnvironment,Int32).0.this\.\_environment\ := \Unum::.ctor(UnumEnvironment,Int32).0.environment\;
                        \Unum::.ctor(UnumEnvironment,Int32).0.array33fbc39d577dad5ed6f3add64bb11d85840cbcf74dc3de0631f99002274571ae\ := (others => to_unsigned(0, 32));
                        \Unum::.ctor(UnumEnvironment,Int32).0.array33fbc39d577dad5ed6f3add64bb11d85840cbcf74dc3de0631f99002274571ae\(to_integer(to_signed(0, 32))) := unsigned(\Unum::.ctor(UnumEnvironment,Int32).0.value\);
                        \Unum::.ctor(UnumEnvironment,Int32).0.arrayc56f74e3798679843c34bc7afcaef2219b75aeedea3562d19b496a830cfa8fe8\ := (others => to_unsigned(0, 32));
                        \Unum::.ctor(UnumEnvironment,Int32).0.arrayc56f74e3798679843c34bc7afcaef2219b75aeedea3562d19b496a830cfa8fe8\(to_integer(to_signed(0, 32))) := unsigned(signed(0 - unsigned(\Unum::.ctor(UnumEnvironment,Int32).0.value\)));
                        \Unum::.ctor(UnumEnvironment,Int32).0.binaryOperationResult.0\ := \Unum::.ctor(UnumEnvironment,Int32).0.value\ >= to_signed(0, 32);

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \Unum::.ctor(UnumEnvironment,Int32).0._State_4\ and ends in state \Unum::.ctor(UnumEnvironment,Int32).0._State_5\.
                        --     * The false branch starts in state \Unum::.ctor(UnumEnvironment,Int32).0._State_6\ and ends in state \Unum::.ctor(UnumEnvironment,Int32).0._State_7\.
                        --     * Execution after either branch will continue in the following state: \Unum::.ctor(UnumEnvironment,Int32).0._State_3\.

                        if (\Unum::.ctor(UnumEnvironment,Int32).0.binaryOperationResult.0\) then 
                            \Unum::.ctor(UnumEnvironment,Int32).0._State\ := \Unum::.ctor(UnumEnvironment,Int32).0._State_4\;
                        else 
                            \Unum::.ctor(UnumEnvironment,Int32).0._State\ := \Unum::.ctor(UnumEnvironment,Int32).0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \Unum::.ctor(UnumEnvironment,Int32).0._State_3\ => 
                        -- State after the if-else which was started in state \Unum::.ctor(UnumEnvironment,Int32).0._State_2\.
                        \Unum::.ctor(UnumEnvironment,Int32).0.this\.\UnumBits\ := \Unum::.ctor(UnumEnvironment,Int32).0.conditional65ed64d003b02a249ce90498ecf1a8ab72b84c723e77e357f582c5a48bb18fc1\;
                        \Unum::.ctor(UnumEnvironment,Int32).0._State\ := \Unum::.ctor(UnumEnvironment,Int32).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,Int32).0._State_4\ => 
                        -- True branch of the if-else started in state \Unum::.ctor(UnumEnvironment,Int32).0._State_2\.
                        -- Initializing record fields to their defaults.
                        \Unum::.ctor(UnumEnvironment,Int32).0.object739e7c0ee2e2d7e2885cba3d8567c7f7fc002803beba2f5f98ae4af41e10ce82\.\IsNull\ := false;
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.UInt32[],System.Boolean)
                        \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).this.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,Int32).0.object739e7c0ee2e2d7e2885cba3d8567c7f7fc002803beba2f5f98ae4af41e10ce82\;
                        \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).environment.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,Int32).0.environment\;
                        \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).value.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,Int32).0.array33fbc39d577dad5ed6f3add64bb11d85840cbcf74dc3de0631f99002274571ae\;
                        \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).negative.parameter.Out.0\ <= False;
                        \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean)._Started.0\ <= true;
                        \Unum::.ctor(UnumEnvironment,Int32).0._State\ := \Unum::.ctor(UnumEnvironment,Int32).0._State_5\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,Int32).0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.UInt32[],System.Boolean)
                        if (\Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean)._Started.0\ = \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean)._Finished.0\) then 
                            \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean)._Started.0\ <= false;
                            \Unum::.ctor(UnumEnvironment,Int32).0.object739e7c0ee2e2d7e2885cba3d8567c7f7fc002803beba2f5f98ae4af41e10ce82\ := \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).this.parameter.In.0\;
                            \Unum::.ctor(UnumEnvironment,Int32).0.environment\ := \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).environment.parameter.In.0\;
                            \Unum::.ctor(UnumEnvironment,Int32).0.array33fbc39d577dad5ed6f3add64bb11d85840cbcf74dc3de0631f99002274571ae\ := \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).value.parameter.In.0\;
                            \Unum::.ctor(UnumEnvironment,Int32).0.conditional65ed64d003b02a249ce90498ecf1a8ab72b84c723e77e357f582c5a48bb18fc1\ := \Unum::.ctor(UnumEnvironment,Int32).0.object739e7c0ee2e2d7e2885cba3d8567c7f7fc002803beba2f5f98ae4af41e10ce82\.\UnumBits\;
                            -- Going to the state after the if-else which was started in state \Unum::.ctor(UnumEnvironment,Int32).0._State_2\.
                            if (\Unum::.ctor(UnumEnvironment,Int32).0._State\ = \Unum::.ctor(UnumEnvironment,Int32).0._State_5\) then 
                                \Unum::.ctor(UnumEnvironment,Int32).0._State\ := \Unum::.ctor(UnumEnvironment,Int32).0._State_3\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,Int32).0._State_6\ => 
                        -- False branch of the if-else started in state \Unum::.ctor(UnumEnvironment,Int32).0._State_2\.
                        -- Initializing record fields to their defaults.
                        \Unum::.ctor(UnumEnvironment,Int32).0.object308d6421e1cd9a8ca8e86fd94126f7dddd720821b3965d0d437be91e799be3b9\.\IsNull\ := false;
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.UInt32[],System.Boolean)
                        \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).this.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,Int32).0.object308d6421e1cd9a8ca8e86fd94126f7dddd720821b3965d0d437be91e799be3b9\;
                        \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).environment.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,Int32).0.environment\;
                        \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).value.parameter.Out.0\ <= \Unum::.ctor(UnumEnvironment,Int32).0.arrayc56f74e3798679843c34bc7afcaef2219b75aeedea3562d19b496a830cfa8fe8\;
                        \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).negative.parameter.Out.0\ <= True;
                        \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean)._Started.0\ <= true;
                        \Unum::.ctor(UnumEnvironment,Int32).0._State\ := \Unum::.ctor(UnumEnvironment,Int32).0._State_7\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::.ctor(UnumEnvironment,Int32).0._State_7\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.UInt32[],System.Boolean)
                        if (\Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean)._Started.0\ = \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean)._Finished.0\) then 
                            \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean)._Started.0\ <= false;
                            \Unum::.ctor(UnumEnvironment,Int32).0.object308d6421e1cd9a8ca8e86fd94126f7dddd720821b3965d0d437be91e799be3b9\ := \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).this.parameter.In.0\;
                            \Unum::.ctor(UnumEnvironment,Int32).0.environment\ := \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).environment.parameter.In.0\;
                            \Unum::.ctor(UnumEnvironment,Int32).0.arrayc56f74e3798679843c34bc7afcaef2219b75aeedea3562d19b496a830cfa8fe8\ := \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).value.parameter.In.0\;
                            \Unum::.ctor(UnumEnvironment,Int32).0.conditional65ed64d003b02a249ce90498ecf1a8ab72b84c723e77e357f582c5a48bb18fc1\ := \Unum::.ctor(UnumEnvironment,Int32).0.object308d6421e1cd9a8ca8e86fd94126f7dddd720821b3965d0d437be91e799be3b9\.\UnumBits\;
                            -- Going to the state after the if-else which was started in state \Unum::.ctor(UnumEnvironment,Int32).0._State_2\.
                            if (\Unum::.ctor(UnumEnvironment,Int32).0._State\ = \Unum::.ctor(UnumEnvironment,Int32).0._State_7\) then 
                                \Unum::.ctor(UnumEnvironment,Int32).0._State\ := \Unum::.ctor(UnumEnvironment,Int32).0._State_3\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.Int32).0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::SetUnumBits(System.Boolean,Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean,System.Byte,System.UInt16).0 state machine start
    \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._StateMachine\: process (\Clock\) 
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\: \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._States\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_0\;
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.this\: \Lombiq.Unum.Unum\;
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.signBit\: boolean := false;
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.exponent\: \Lombiq.Unum.BitMask\;
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.fraction\: \Lombiq.Unum.BitMask\;
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.uncertainityBit\: boolean := false;
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.exponentSize\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.fractionSize\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.bitMask\: \Lombiq.Unum.BitMask\;
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.array8756220799ceaafd5b50dac1ff26f31915dcc57cd912ca3e7d8bfd1b17d2f16e\: \unsigned32_Array\(0 to 0) := (others => to_unsigned(0, 32));
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.object3efd49a19499cd5d8cc4aa1d852393f30b746e0ccd1de8def3509997f3c7f683\: \Lombiq.Unum.BitMask\;
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.1\: \Lombiq.Unum.BitMask\;
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.2\: \Lombiq.Unum.BitMask\;
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.3\: \Lombiq.Unum.BitMask\;
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.4\: \Lombiq.Unum.BitMask\;
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.5\: \Lombiq.Unum.BitMask\;
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.6\: \Lombiq.Unum.BitMask\;
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.binaryOperationResult.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.binaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.7\: \Lombiq.Unum.BitMask\;
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.8\: \Lombiq.Unum.BitMask\;
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.9\: \Lombiq.Unum.BitMask\;
        Variable \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.10\: \Lombiq.Unum.BitMask\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._Finished\ <= false;
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_Size()._Started.0\ <= false;
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 32));
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\ <= to_signed(0, 32);
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= false;
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\ <= to_unsigned(0, 32);
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ <= false;
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_UncertaintyBitMask()._Started.0\ <= false;
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= false;
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_SignBitMask()._Started.0\ <= false;
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_0\;
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.signBit\ := false;
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.uncertainityBit\ := false;
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.exponentSize\ := to_unsigned(0, 8);
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.fractionSize\ := to_unsigned(0, 16);
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.array8756220799ceaafd5b50dac1ff26f31915dcc57cd912ca3e7d8bfd1b17d2f16e\ := (others => to_unsigned(0, 32));
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.0\ := to_unsigned(0, 16);
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.binaryOperationResult.0\ := to_unsigned(0, 16);
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.binaryOperationResult.1\ := to_signed(0, 32);
            else 
                case \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ is 
                    when \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._Started\ = true) then 
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._Started\ = true) then 
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._Finished\ <= true;
                        else 
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._Finished\ <= false;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_2\ => 
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.this\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.this.parameter.In\;
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.signBit\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.signBit.parameter.In\;
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.exponent\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.exponent.parameter.In\;
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.fraction\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.fraction.parameter.In\;
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.uncertainityBit\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.uncertainityBit.parameter.In\;
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.exponentSize\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.exponentSize.parameter.In\;
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.fractionSize\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.fractionSize.parameter.In\;
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.array8756220799ceaafd5b50dac1ff26f31915dcc57cd912ca3e7d8bfd1b17d2f16e\ := (others => to_unsigned(0, 32));
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.array8756220799ceaafd5b50dac1ff26f31915dcc57cd912ca3e7d8bfd1b17d2f16e\(to_integer(to_signed(0, 32))) := resize(\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.exponentSize\, 32);
                        -- Initializing record fields to their defaults.
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.object3efd49a19499cd5d8cc4aa1d852393f30b746e0ccd1de8def3509997f3c7f683\.\IsNull\ := false;
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.object3efd49a19499cd5d8cc4aa1d852393f30b746e0ccd1de8def3509997f3c7f683\.\Size\ := to_unsigned(0, 16);
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.object3efd49a19499cd5d8cc4aa1d852393f30b746e0ccd1de8def3509997f3c7f683\.\SegmentCount\ := to_unsigned(0, 16);
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.object3efd49a19499cd5d8cc4aa1d852393f30b746e0ccd1de8def3509997f3c7f683\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::get_Size()
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_Size().this.parameter.Out.0\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.this\;
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_Size()._Started.0\ <= true;
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::get_Size()
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_Size()._Started.0\ = \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_Size()._Finished.0\) then 
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_Size()._Started.0\ <= false;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.0\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_Size().return.0\;
                            -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.object3efd49a19499cd5d8cc4aa1d852393f30b746e0ccd1de8def3509997f3c7f683\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\(0 to 0) <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.array8756220799ceaafd5b50dac1ff26f31915dcc57cd912ca3e7d8bfd1b17d2f16e\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.0\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= true;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\) then 
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.object3efd49a19499cd5d8cc4aa1d852393f30b746e0ccd1de8def3509997f3c7f683\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.array8756220799ceaafd5b50dac1ff26f31915dcc57cd912ca3e7d8bfd1b17d2f16e\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\(0 to 0);
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.object3efd49a19499cd5d8cc4aa1d852393f30b746e0ccd1de8def3509997f3c7f683\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\ <= to_signed(8, 32);
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= true;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ = \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\) then 
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= false;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.1\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32).return.0\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.bitMask\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.1\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,System.UInt32)
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,UInt32).left.parameter.Out.0\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.bitMask\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\ <= resize(\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.fractionSize\, 32);
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ <= true;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_6\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,System.UInt32)
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ = \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\) then 
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ <= false;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.2\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,UInt32).return.0\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.bitMask\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.2\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_8\ and ends in state \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_10\.
                            --     * Execution after either branch will continue in the following state: \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_7\.

                            if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.uncertainityBit\) then 
                                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_8\;
                            else 
                                -- There was no false branch, so going directly to the state after the if-else.
                                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_7\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_7\ => 
                        -- State after the if-else which was started in state \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_6\.
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.fraction\;
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\ <= to_signed(13, 32);
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= true;
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_11\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_8\ => 
                        -- True branch of the if-else started in state \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_6\.
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_UncertaintyBitMask()
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_UncertaintyBitMask().this.parameter.Out.0\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.this\;
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_UncertaintyBitMask()._Started.0\ <= true;
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_9\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_9\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_UncertaintyBitMask()
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_UncertaintyBitMask()._Started.0\ = \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_UncertaintyBitMask()._Finished.0\) then 
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_UncertaintyBitMask()._Started.0\ <= false;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.3\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_UncertaintyBitMask().return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask).left.parameter.Out.0\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.bitMask\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask).right.parameter.Out.0\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.3\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= true;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_10\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_10\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ = \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\) then 
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= false;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.4\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask).return.0\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.bitMask\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.4\;
                            -- Going to the state after the if-else which was started in state \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_6\.
                            if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ = \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_10\) then 
                                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_7\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_11\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ = \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\) then 
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= false;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.5\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32).return.0\;
                            -- The last invocation for the target state machine finished in the previous state, so need to start the next one in the next state.
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_12\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_12\ => 
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask).left.parameter.Out.0\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.bitMask\;
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask).right.parameter.Out.0\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.5\;
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= true;
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_13\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_13\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ = \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\) then 
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= false;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.6\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask).return.0\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.bitMask\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.6\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.binaryOperationResult.0\ := to_unsigned(13, 16) + \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.fractionSize\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.binaryOperationResult.1\ := resize(signed(\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.binaryOperationResult.0\ + to_unsigned(1, 16)), 32);
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.exponent\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\ <= (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.binaryOperationResult.1\);
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= true;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_14\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_14\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ = \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\) then 
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= false;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.7\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32).return.0\;
                            -- The last invocation for the target state machine finished in the previous state, so need to start the next one in the next state.
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_15\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_15\ => 
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask).left.parameter.Out.0\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.bitMask\;
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask).right.parameter.Out.0\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.7\;
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= true;
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_16\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_16\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ = \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\) then 
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= false;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.8\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask).return.0\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.bitMask\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.8\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_18\ and ends in state \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_20\.
                            --     * Execution after either branch will continue in the following state: \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_17\.

                            if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.signBit\) then 
                                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_18\;
                            else 
                                -- There was no false branch, so going directly to the state after the if-else.
                                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_17\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_17\ => 
                        -- State after the if-else which was started in state \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_16\.
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.bitMask\;
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_18\ => 
                        -- True branch of the if-else started in state \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_16\.
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_SignBitMask()
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_SignBitMask().this.parameter.Out.0\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.this\;
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_SignBitMask()._Started.0\ <= true;
                        \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_19\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_19\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_SignBitMask()
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_SignBitMask()._Started.0\ = \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_SignBitMask()._Finished.0\) then 
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_SignBitMask()._Started.0\ <= false;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.9\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_SignBitMask().return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask).left.parameter.Out.0\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.bitMask\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask).right.parameter.Out.0\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.9\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= true;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_20\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_20\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ = \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\) then 
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= false;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.10\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask).return.0\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.bitMask\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return.10\;
                            -- Going to the state after the if-else which was started in state \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_16\.
                            if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ = \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_20\) then 
                                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State\ := \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._State_17\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::SetUnumBits(System.Boolean,Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean,System.Byte,System.UInt16).0 state machine end


    -- System.UInt32[] Lombiq.Unum.Unum::FractionToUintArray().0 state machine start
    \Unum::FractionToUintArray().0._StateMachine\: process (\Clock\) 
        Variable \Unum::FractionToUintArray().0._State\: \Unum::FractionToUintArray().0._States\ := \Unum::FractionToUintArray().0._State_0\;
        Variable \Unum::FractionToUintArray().0.this\: \Lombiq.Unum.Unum\;
        Variable \Unum::FractionToUintArray().0.bitMask\: \Lombiq.Unum.BitMask\;
        Variable \Unum::FractionToUintArray().0.array\: \unsigned32_Array\(0 to 8) := (others => to_unsigned(0, 32));
        Variable \Unum::FractionToUintArray().0.i\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::FractionToUintArray().0.flag\: boolean := false;
        Variable \Unum::FractionToUintArray().0.return.0\: \Lombiq.Unum.BitMask\;
        Variable \Unum::FractionToUintArray().0.return.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::FractionToUintArray().0.return.2\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::FractionToUintArray().0.binaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::FractionToUintArray().0.return.3\: \Lombiq.Unum.BitMask\;
        Variable \Unum::FractionToUintArray().0.binaryOperationResult.1\: boolean := false;
        Variable \Unum::FractionToUintArray().0.binaryOperationResult.2\: boolean := false;
        Variable \Unum::FractionToUintArray().0.binaryOperationResult.3\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::FractionToUintArray().0.return.4\: boolean := false;
        Variable \Unum::FractionToUintArray().0.binaryOperationResult.4\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::FractionToUintArray().0.binaryOperationResult.5\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::FractionToUintArray().0.binaryOperationResult.6\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Unum::FractionToUintArray().0.binaryOperationResult.7\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::FractionToUintArray().0.binaryOperationResult.8\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::FractionToUintArray().0.binaryOperationResult.9\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Unum::FractionToUintArray().0.binaryOperationResult.10\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::FractionToUintArray().0.binaryOperationResult.11\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::FractionToUintArray().0.binaryOperationResult.12\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::FractionToUintArray().0._Finished\ <= false;
                \Unum::FractionToUintArray().0.return\ <= (others => to_unsigned(0, 32));
                \Unum::FractionToUintArray().0.Unum::FractionWithHiddenBit()._Started.0\ <= false;
                \Unum::FractionToUintArray().0.Unum::ExponentValueWithBias()._Started.0\ <= false;
                \Unum::FractionToUintArray().0.Unum::FractionSize()._Started.0\ <= false;
                \Unum::FractionToUintArray().0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\ <= to_signed(0, 32);
                \Unum::FractionToUintArray().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= false;
                \Unum::FractionToUintArray().0.Unum::IsPositive()._Started.0\ <= false;
                \Unum::FractionToUintArray().0._State\ := \Unum::FractionToUintArray().0._State_0\;
                \Unum::FractionToUintArray().0.array\ := (others => to_unsigned(0, 32));
                \Unum::FractionToUintArray().0.i\ := to_signed(0, 32);
                \Unum::FractionToUintArray().0.flag\ := false;
                \Unum::FractionToUintArray().0.return.1\ := to_signed(0, 32);
                \Unum::FractionToUintArray().0.return.2\ := to_unsigned(0, 16);
                \Unum::FractionToUintArray().0.binaryOperationResult.0\ := to_signed(0, 32);
                \Unum::FractionToUintArray().0.binaryOperationResult.1\ := false;
                \Unum::FractionToUintArray().0.binaryOperationResult.2\ := false;
                \Unum::FractionToUintArray().0.binaryOperationResult.3\ := to_signed(0, 32);
                \Unum::FractionToUintArray().0.return.4\ := false;
                \Unum::FractionToUintArray().0.binaryOperationResult.4\ := to_signed(0, 32);
                \Unum::FractionToUintArray().0.binaryOperationResult.5\ := to_signed(0, 32);
                \Unum::FractionToUintArray().0.binaryOperationResult.6\ := to_unsigned(0, 32);
                \Unum::FractionToUintArray().0.binaryOperationResult.7\ := to_signed(0, 32);
                \Unum::FractionToUintArray().0.binaryOperationResult.8\ := to_signed(0, 32);
                \Unum::FractionToUintArray().0.binaryOperationResult.9\ := to_unsigned(0, 32);
                \Unum::FractionToUintArray().0.binaryOperationResult.10\ := to_signed(0, 32);
                \Unum::FractionToUintArray().0.binaryOperationResult.11\ := to_signed(0, 32);
                \Unum::FractionToUintArray().0.binaryOperationResult.12\ := to_unsigned(0, 32);
            else 
                case \Unum::FractionToUintArray().0._State\ is 
                    when \Unum::FractionToUintArray().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::FractionToUintArray().0._Started\ = true) then 
                            \Unum::FractionToUintArray().0._State\ := \Unum::FractionToUintArray().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionToUintArray().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::FractionToUintArray().0._Started\ = true) then 
                            \Unum::FractionToUintArray().0._Finished\ <= true;
                        else 
                            \Unum::FractionToUintArray().0._Finished\ <= false;
                            \Unum::FractionToUintArray().0._State\ := \Unum::FractionToUintArray().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionToUintArray().0._State_2\ => 
                        \Unum::FractionToUintArray().0.this\ := \Unum::FractionToUintArray().0.this.parameter.In\;
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit()
                        \Unum::FractionToUintArray().0.Unum::FractionWithHiddenBit().this.parameter.Out.0\ <= \Unum::FractionToUintArray().0.this\;
                        \Unum::FractionToUintArray().0.Unum::FractionWithHiddenBit()._Started.0\ <= true;
                        \Unum::FractionToUintArray().0._State\ := \Unum::FractionToUintArray().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionToUintArray().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit()
                        if (\Unum::FractionToUintArray().0.Unum::FractionWithHiddenBit()._Started.0\ = \Unum::FractionToUintArray().0.Unum::FractionWithHiddenBit()._Finished.0\) then 
                            \Unum::FractionToUintArray().0.Unum::FractionWithHiddenBit()._Started.0\ <= false;
                            \Unum::FractionToUintArray().0.return.0\ := \Unum::FractionToUintArray().0.Unum::FractionWithHiddenBit().return.0\;
                            -- Starting state machine invocation for the following method: System.Int32 Lombiq.Unum.Unum::ExponentValueWithBias()
                            \Unum::FractionToUintArray().0.Unum::ExponentValueWithBias().this.parameter.Out.0\ <= \Unum::FractionToUintArray().0.this\;
                            \Unum::FractionToUintArray().0.Unum::ExponentValueWithBias()._Started.0\ <= true;
                            \Unum::FractionToUintArray().0._State\ := \Unum::FractionToUintArray().0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionToUintArray().0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Int32 Lombiq.Unum.Unum::ExponentValueWithBias()
                        if (\Unum::FractionToUintArray().0.Unum::ExponentValueWithBias()._Started.0\ = \Unum::FractionToUintArray().0.Unum::ExponentValueWithBias()._Finished.0\) then 
                            \Unum::FractionToUintArray().0.Unum::ExponentValueWithBias()._Started.0\ <= false;
                            \Unum::FractionToUintArray().0.return.1\ := \Unum::FractionToUintArray().0.Unum::ExponentValueWithBias().return.0\;
                            -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::FractionSize()
                            \Unum::FractionToUintArray().0.Unum::FractionSize().this.parameter.Out.0\ <= \Unum::FractionToUintArray().0.this\;
                            \Unum::FractionToUintArray().0.Unum::FractionSize()._Started.0\ <= true;
                            \Unum::FractionToUintArray().0._State\ := \Unum::FractionToUintArray().0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionToUintArray().0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::FractionSize()
                        if (\Unum::FractionToUintArray().0.Unum::FractionSize()._Started.0\ = \Unum::FractionToUintArray().0.Unum::FractionSize()._Finished.0\) then 
                            \Unum::FractionToUintArray().0.Unum::FractionSize()._Started.0\ <= false;
                            \Unum::FractionToUintArray().0.return.2\ := \Unum::FractionToUintArray().0.Unum::FractionSize().return.0\;
                            \Unum::FractionToUintArray().0.binaryOperationResult.0\ := resize(\Unum::FractionToUintArray().0.return.1\ - resize(signed(\Unum::FractionToUintArray().0.return.2\), 32), 32);
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                            \Unum::FractionToUintArray().0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\ <= \Unum::FractionToUintArray().0.return.0\;
                            \Unum::FractionToUintArray().0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\ <= \Unum::FractionToUintArray().0.binaryOperationResult.0\;
                            \Unum::FractionToUintArray().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= true;
                            \Unum::FractionToUintArray().0._State\ := \Unum::FractionToUintArray().0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::FractionToUintArray().0._State_6\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                        if (\Unum::FractionToUintArray().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ = \Unum::FractionToUintArray().0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\) then 
                            \Unum::FractionToUintArray().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= false;
                            \Unum::FractionToUintArray().0.return.3\ := \Unum::FractionToUintArray().0.BitMask::op_LeftShift(BitMask,Int32).return.0\;
                            \Unum::FractionToUintArray().0.bitMask\ := \Unum::FractionToUintArray().0.return.3\;
                            \Unum::FractionToUintArray().0.array\ := (others => to_unsigned(0, 32));
                            \Unum::FractionToUintArray().0.i\ := to_signed(0, 32);
                            -- Starting a while loop.
                            -- The while loop's condition (also added here to be able to branch off early if the loop body shouldn't be executed at all):
                            \Unum::FractionToUintArray().0.binaryOperationResult.1\ := \Unum::FractionToUintArray().0.i\ < resize(signed(\Unum::FractionToUintArray().0.bitMask\.\SegmentCount\), 32);
                            if (\Unum::FractionToUintArray().0.binaryOperationResult.1\) then 
                                \Unum::FractionToUintArray().0._State\ := \Unum::FractionToUintArray().0._State_7\;
                            else 
                                \Unum::FractionToUintArray().0._State\ := \Unum::FractionToUintArray().0._State_8\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::FractionToUintArray().0._State_7\ => 
                        -- Repeated state of the while loop which was started in state \Unum::FractionToUintArray().0._State_6\.
                        -- The while loop's condition:
                        \Unum::FractionToUintArray().0.binaryOperationResult.2\ := \Unum::FractionToUintArray().0.i\ < resize(signed(\Unum::FractionToUintArray().0.bitMask\.\SegmentCount\), 32);
                        if (\Unum::FractionToUintArray().0.binaryOperationResult.2\) then 
                            \Unum::FractionToUintArray().0.array\(to_integer(\Unum::FractionToUintArray().0.i\)) := \Unum::FractionToUintArray().0.bitMask\.\Segments\(to_integer(\Unum::FractionToUintArray().0.i\));
                            \Unum::FractionToUintArray().0.binaryOperationResult.3\ := \Unum::FractionToUintArray().0.i\ + to_signed(1, 32);
                            \Unum::FractionToUintArray().0.i\ := \Unum::FractionToUintArray().0.binaryOperationResult.3\;
                        else 
                            \Unum::FractionToUintArray().0._State\ := \Unum::FractionToUintArray().0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \Unum::FractionToUintArray().0._State_8\ => 
                        -- State after the while loop which was started in state \Unum::FractionToUintArray().0._State_6\.
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::IsPositive()
                        \Unum::FractionToUintArray().0.Unum::IsPositive().this.parameter.Out.0\ <= \Unum::FractionToUintArray().0.this\;
                        \Unum::FractionToUintArray().0.Unum::IsPositive()._Started.0\ <= true;
                        \Unum::FractionToUintArray().0._State\ := \Unum::FractionToUintArray().0._State_9\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::FractionToUintArray().0._State_9\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::IsPositive()
                        if (\Unum::FractionToUintArray().0.Unum::IsPositive()._Started.0\ = \Unum::FractionToUintArray().0.Unum::IsPositive()._Finished.0\) then 
                            \Unum::FractionToUintArray().0.Unum::IsPositive()._Started.0\ <= false;
                            \Unum::FractionToUintArray().0.return.4\ := \Unum::FractionToUintArray().0.Unum::IsPositive().return.0\;
                            \Unum::FractionToUintArray().0.flag\ := not(\Unum::FractionToUintArray().0.return.4\);

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::FractionToUintArray().0._State_11\ and ends in state \Unum::FractionToUintArray().0._State_11\.
                            --     * The false branch starts in state \Unum::FractionToUintArray().0._State_12\ and ends in state \Unum::FractionToUintArray().0._State_12\.
                            --     * Execution after either branch will continue in the following state: \Unum::FractionToUintArray().0._State_10\.

                            if (\Unum::FractionToUintArray().0.flag\) then 
                                \Unum::FractionToUintArray().0._State\ := \Unum::FractionToUintArray().0._State_11\;
                            else 
                                \Unum::FractionToUintArray().0._State\ := \Unum::FractionToUintArray().0._State_12\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionToUintArray().0._State_10\ => 
                        -- State after the if-else which was started in state \Unum::FractionToUintArray().0._State_9\.
                        \Unum::FractionToUintArray().0.return\ <= \Unum::FractionToUintArray().0.array\;
                        \Unum::FractionToUintArray().0._State\ := \Unum::FractionToUintArray().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionToUintArray().0._State_11\ => 
                        -- True branch of the if-else started in state \Unum::FractionToUintArray().0._State_9\.
                        \Unum::FractionToUintArray().0.binaryOperationResult.4\ := resize(signed(\Unum::FractionToUintArray().0.bitMask\.\SegmentCount\ - to_unsigned(1, 16)), 32);
                        \Unum::FractionToUintArray().0.binaryOperationResult.5\ := resize(signed(\Unum::FractionToUintArray().0.bitMask\.\SegmentCount\ - to_unsigned(1, 16)), 32);
                        -- Since the integer literal 2147483648 was out of the VHDL integer range it was substituted with a binary literal (10000000000000000000000000000000).
                        \Unum::FractionToUintArray().0.binaryOperationResult.6\ := \Unum::FractionToUintArray().0.array\(to_integer((\Unum::FractionToUintArray().0.binaryOperationResult.5\))) or "10000000000000000000000000000000";
                        \Unum::FractionToUintArray().0.array\(to_integer((\Unum::FractionToUintArray().0.binaryOperationResult.4\))) := \Unum::FractionToUintArray().0.binaryOperationResult.6\;
                        -- Going to the state after the if-else which was started in state \Unum::FractionToUintArray().0._State_9\.
                        if (\Unum::FractionToUintArray().0._State\ = \Unum::FractionToUintArray().0._State_11\) then 
                            \Unum::FractionToUintArray().0._State\ := \Unum::FractionToUintArray().0._State_10\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \Unum::FractionToUintArray().0._State_12\ => 
                        -- False branch of the if-else started in state \Unum::FractionToUintArray().0._State_9\.
                        \Unum::FractionToUintArray().0.binaryOperationResult.7\ := resize(signed(\Unum::FractionToUintArray().0.bitMask\.\SegmentCount\ - to_unsigned(1, 16)), 32);
                        \Unum::FractionToUintArray().0.binaryOperationResult.8\ := resize(signed(\Unum::FractionToUintArray().0.bitMask\.\SegmentCount\ - to_unsigned(1, 16)), 32);
                        \Unum::FractionToUintArray().0.binaryOperationResult.9\ := shift_left(\Unum::FractionToUintArray().0.array\(to_integer((\Unum::FractionToUintArray().0.binaryOperationResult.8\))), to_integer(to_signed(1, 32)));
                        \Unum::FractionToUintArray().0.array\(to_integer((\Unum::FractionToUintArray().0.binaryOperationResult.7\))) := \Unum::FractionToUintArray().0.binaryOperationResult.9\;
                        \Unum::FractionToUintArray().0.binaryOperationResult.10\ := resize(signed(\Unum::FractionToUintArray().0.bitMask\.\SegmentCount\ - to_unsigned(1, 16)), 32);
                        \Unum::FractionToUintArray().0.binaryOperationResult.11\ := resize(signed(\Unum::FractionToUintArray().0.bitMask\.\SegmentCount\ - to_unsigned(1, 16)), 32);
                        \Unum::FractionToUintArray().0.binaryOperationResult.12\ := shift_right(\Unum::FractionToUintArray().0.array\(to_integer((\Unum::FractionToUintArray().0.binaryOperationResult.11\))), to_integer(to_signed(1, 32)));
                        \Unum::FractionToUintArray().0.array\(to_integer((\Unum::FractionToUintArray().0.binaryOperationResult.10\))) := \Unum::FractionToUintArray().0.binaryOperationResult.12\;
                        -- Going to the state after the if-else which was started in state \Unum::FractionToUintArray().0._State_9\.
                        if (\Unum::FractionToUintArray().0._State\ = \Unum::FractionToUintArray().0._State_12\) then 
                            \Unum::FractionToUintArray().0._State\ := \Unum::FractionToUintArray().0._State_10\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.6
                end case;
            end if;
        end if;
    end process;
    -- System.UInt32[] Lombiq.Unum.Unum::FractionToUintArray().0 state machine end


    -- System.Boolean Lombiq.Unum.Unum::IsExact().0 state machine start
    \Unum::IsExact().0._StateMachine\: process (\Clock\) 
        Variable \Unum::IsExact().0._State\: \Unum::IsExact().0._States\ := \Unum::IsExact().0._State_0\;
        Variable \Unum::IsExact().0.this\: \Lombiq.Unum.Unum\;
        Variable \Unum::IsExact().0.return.0\: \Lombiq.Unum.BitMask\;
        Variable \Unum::IsExact().0.return.1\: \Lombiq.Unum.BitMask\;
        Variable \Unum::IsExact().0.return.2\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::IsExact().0._Finished\ <= false;
                \Unum::IsExact().0.return\ <= false;
                \Unum::IsExact().0.Unum::get_UncertaintyBitMask()._Started.0\ <= false;
                \Unum::IsExact().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ <= false;
                \Unum::IsExact().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ <= false;
                \Unum::IsExact().0._State\ := \Unum::IsExact().0._State_0\;
                \Unum::IsExact().0.return.2\ := false;
            else 
                case \Unum::IsExact().0._State\ is 
                    when \Unum::IsExact().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::IsExact().0._Started\ = true) then 
                            \Unum::IsExact().0._State\ := \Unum::IsExact().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsExact().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::IsExact().0._Started\ = true) then 
                            \Unum::IsExact().0._Finished\ <= true;
                        else 
                            \Unum::IsExact().0._Finished\ <= false;
                            \Unum::IsExact().0._State\ := \Unum::IsExact().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsExact().0._State_2\ => 
                        \Unum::IsExact().0.this\ := \Unum::IsExact().0.this.parameter.In\;
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_UncertaintyBitMask()
                        \Unum::IsExact().0.Unum::get_UncertaintyBitMask().this.parameter.Out.0\ <= \Unum::IsExact().0.this\;
                        \Unum::IsExact().0.Unum::get_UncertaintyBitMask()._Started.0\ <= true;
                        \Unum::IsExact().0._State\ := \Unum::IsExact().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsExact().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_UncertaintyBitMask()
                        if (\Unum::IsExact().0.Unum::get_UncertaintyBitMask()._Started.0\ = \Unum::IsExact().0.Unum::get_UncertaintyBitMask()._Finished.0\) then 
                            \Unum::IsExact().0.Unum::get_UncertaintyBitMask()._Started.0\ <= false;
                            \Unum::IsExact().0.return.0\ := \Unum::IsExact().0.Unum::get_UncertaintyBitMask().return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseAnd(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \Unum::IsExact().0.BitMask::op_BitwiseAnd(BitMask,BitMask).left.parameter.Out.0\ <= \Unum::IsExact().0.this\.\UnumBits\;
                            \Unum::IsExact().0.BitMask::op_BitwiseAnd(BitMask,BitMask).right.parameter.Out.0\ <= \Unum::IsExact().0.return.0\;
                            \Unum::IsExact().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ <= true;
                            \Unum::IsExact().0._State\ := \Unum::IsExact().0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsExact().0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseAnd(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\Unum::IsExact().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ = \Unum::IsExact().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\) then 
                            \Unum::IsExact().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ <= false;
                            \Unum::IsExact().0.return.1\ := \Unum::IsExact().0.BitMask::op_BitwiseAnd(BitMask,BitMask).return.0\;
                            -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.BitMask::op_Equality(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \Unum::IsExact().0.BitMask::op_Equality(BitMask,BitMask).left.parameter.Out.0\ <= \Unum::IsExact().0.return.1\;
                            \Unum::IsExact().0.BitMask::op_Equality(BitMask,BitMask).right.parameter.Out.0\ <= \Unum::IsExact().0.this\.\_environment\.\EmptyBitMask\;
                            \Unum::IsExact().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ <= true;
                            \Unum::IsExact().0._State\ := \Unum::IsExact().0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsExact().0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.BitMask::op_Equality(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\Unum::IsExact().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ = \Unum::IsExact().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\) then 
                            \Unum::IsExact().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ <= false;
                            \Unum::IsExact().0.return.2\ := \Unum::IsExact().0.BitMask::op_Equality(BitMask,BitMask).return.0\;
                            \Unum::IsExact().0.return\ <= \Unum::IsExact().0.return.2\;
                            \Unum::IsExact().0._State\ := \Unum::IsExact().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Lombiq.Unum.Unum::IsExact().0 state machine end


    -- System.Boolean Lombiq.Unum.Unum::IsPositive().0 state machine start
    \Unum::IsPositive().0._StateMachine\: process (\Clock\) 
        Variable \Unum::IsPositive().0._State\: \Unum::IsPositive().0._States\ := \Unum::IsPositive().0._State_0\;
        Variable \Unum::IsPositive().0.this\: \Lombiq.Unum.Unum\;
        Variable \Unum::IsPositive().0.return.0\: \Lombiq.Unum.BitMask\;
        Variable \Unum::IsPositive().0.return.1\: \Lombiq.Unum.BitMask\;
        Variable \Unum::IsPositive().0.return.2\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::IsPositive().0._Finished\ <= false;
                \Unum::IsPositive().0.return\ <= false;
                \Unum::IsPositive().0.Unum::get_SignBitMask()._Started.0\ <= false;
                \Unum::IsPositive().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ <= false;
                \Unum::IsPositive().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ <= false;
                \Unum::IsPositive().0._State\ := \Unum::IsPositive().0._State_0\;
                \Unum::IsPositive().0.return.2\ := false;
            else 
                case \Unum::IsPositive().0._State\ is 
                    when \Unum::IsPositive().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::IsPositive().0._Started\ = true) then 
                            \Unum::IsPositive().0._State\ := \Unum::IsPositive().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsPositive().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::IsPositive().0._Started\ = true) then 
                            \Unum::IsPositive().0._Finished\ <= true;
                        else 
                            \Unum::IsPositive().0._Finished\ <= false;
                            \Unum::IsPositive().0._State\ := \Unum::IsPositive().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsPositive().0._State_2\ => 
                        \Unum::IsPositive().0.this\ := \Unum::IsPositive().0.this.parameter.In\;
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_SignBitMask()
                        \Unum::IsPositive().0.Unum::get_SignBitMask().this.parameter.Out.0\ <= \Unum::IsPositive().0.this\;
                        \Unum::IsPositive().0.Unum::get_SignBitMask()._Started.0\ <= true;
                        \Unum::IsPositive().0._State\ := \Unum::IsPositive().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsPositive().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_SignBitMask()
                        if (\Unum::IsPositive().0.Unum::get_SignBitMask()._Started.0\ = \Unum::IsPositive().0.Unum::get_SignBitMask()._Finished.0\) then 
                            \Unum::IsPositive().0.Unum::get_SignBitMask()._Started.0\ <= false;
                            \Unum::IsPositive().0.return.0\ := \Unum::IsPositive().0.Unum::get_SignBitMask().return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseAnd(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \Unum::IsPositive().0.BitMask::op_BitwiseAnd(BitMask,BitMask).left.parameter.Out.0\ <= \Unum::IsPositive().0.this\.\UnumBits\;
                            \Unum::IsPositive().0.BitMask::op_BitwiseAnd(BitMask,BitMask).right.parameter.Out.0\ <= \Unum::IsPositive().0.return.0\;
                            \Unum::IsPositive().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ <= true;
                            \Unum::IsPositive().0._State\ := \Unum::IsPositive().0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsPositive().0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseAnd(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\Unum::IsPositive().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ = \Unum::IsPositive().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\) then 
                            \Unum::IsPositive().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ <= false;
                            \Unum::IsPositive().0.return.1\ := \Unum::IsPositive().0.BitMask::op_BitwiseAnd(BitMask,BitMask).return.0\;
                            -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.BitMask::op_Equality(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \Unum::IsPositive().0.BitMask::op_Equality(BitMask,BitMask).left.parameter.Out.0\ <= \Unum::IsPositive().0.return.1\;
                            \Unum::IsPositive().0.BitMask::op_Equality(BitMask,BitMask).right.parameter.Out.0\ <= \Unum::IsPositive().0.this\.\_environment\.\EmptyBitMask\;
                            \Unum::IsPositive().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ <= true;
                            \Unum::IsPositive().0._State\ := \Unum::IsPositive().0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsPositive().0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.BitMask::op_Equality(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\Unum::IsPositive().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ = \Unum::IsPositive().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\) then 
                            \Unum::IsPositive().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ <= false;
                            \Unum::IsPositive().0.return.2\ := \Unum::IsPositive().0.BitMask::op_Equality(BitMask,BitMask).return.0\;
                            \Unum::IsPositive().0.return\ <= \Unum::IsPositive().0.return.2\;
                            \Unum::IsPositive().0._State\ := \Unum::IsPositive().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Lombiq.Unum.Unum::IsPositive().0 state machine end


    -- System.Byte Lombiq.Unum.Unum::ExponentSize().0 state machine start
    \Unum::ExponentSize().0._StateMachine\: process (\Clock\) 
        Variable \Unum::ExponentSize().0._State\: \Unum::ExponentSize().0._States\ := \Unum::ExponentSize().0._State_0\;
        Variable \Unum::ExponentSize().0.this\: \Lombiq.Unum.Unum\;
        Variable \Unum::ExponentSize().0.return.0\: \Lombiq.Unum.BitMask\;
        Variable \Unum::ExponentSize().0.return.1\: \Lombiq.Unum.BitMask\;
        Variable \Unum::ExponentSize().0.return.2\: \Lombiq.Unum.BitMask\;
        Variable \Unum::ExponentSize().0.return.3\: \Lombiq.Unum.BitMask\;
        Variable \Unum::ExponentSize().0.return.4\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::ExponentSize().0._Finished\ <= false;
                \Unum::ExponentSize().0.return\ <= to_unsigned(0, 8);
                \Unum::ExponentSize().0.Unum::get_ExponentSizeMask()._Started.0\ <= false;
                \Unum::ExponentSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ <= false;
                \Unum::ExponentSize().0.BitMask::op_RightShift(BitMask,Int32).right.parameter.Out.0\ <= to_signed(0, 32);
                \Unum::ExponentSize().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ <= false;
                \Unum::ExponentSize().0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\ <= to_unsigned(0, 32);
                \Unum::ExponentSize().0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ <= false;
                \Unum::ExponentSize().0.BitMask::GetLowest32Bits()._Started.0\ <= false;
                \Unum::ExponentSize().0._State\ := \Unum::ExponentSize().0._State_0\;
                \Unum::ExponentSize().0.return.4\ := to_unsigned(0, 32);
            else 
                case \Unum::ExponentSize().0._State\ is 
                    when \Unum::ExponentSize().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::ExponentSize().0._Started\ = true) then 
                            \Unum::ExponentSize().0._State\ := \Unum::ExponentSize().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentSize().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::ExponentSize().0._Started\ = true) then 
                            \Unum::ExponentSize().0._Finished\ <= true;
                        else 
                            \Unum::ExponentSize().0._Finished\ <= false;
                            \Unum::ExponentSize().0._State\ := \Unum::ExponentSize().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentSize().0._State_2\ => 
                        \Unum::ExponentSize().0.this\ := \Unum::ExponentSize().0.this.parameter.In\;
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_ExponentSizeMask()
                        \Unum::ExponentSize().0.Unum::get_ExponentSizeMask().this.parameter.Out.0\ <= \Unum::ExponentSize().0.this\;
                        \Unum::ExponentSize().0.Unum::get_ExponentSizeMask()._Started.0\ <= true;
                        \Unum::ExponentSize().0._State\ := \Unum::ExponentSize().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentSize().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_ExponentSizeMask()
                        if (\Unum::ExponentSize().0.Unum::get_ExponentSizeMask()._Started.0\ = \Unum::ExponentSize().0.Unum::get_ExponentSizeMask()._Finished.0\) then 
                            \Unum::ExponentSize().0.Unum::get_ExponentSizeMask()._Started.0\ <= false;
                            \Unum::ExponentSize().0.return.0\ := \Unum::ExponentSize().0.Unum::get_ExponentSizeMask().return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseAnd(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \Unum::ExponentSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask).left.parameter.Out.0\ <= \Unum::ExponentSize().0.this\.\UnumBits\;
                            \Unum::ExponentSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask).right.parameter.Out.0\ <= \Unum::ExponentSize().0.return.0\;
                            \Unum::ExponentSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ <= true;
                            \Unum::ExponentSize().0._State\ := \Unum::ExponentSize().0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentSize().0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseAnd(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\Unum::ExponentSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ = \Unum::ExponentSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\) then 
                            \Unum::ExponentSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ <= false;
                            \Unum::ExponentSize().0.return.1\ := \Unum::ExponentSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask).return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_RightShift(Lombiq.Unum.BitMask,System.Int32)
                            \Unum::ExponentSize().0.BitMask::op_RightShift(BitMask,Int32).left.parameter.Out.0\ <= \Unum::ExponentSize().0.return.1\;
                            \Unum::ExponentSize().0.BitMask::op_RightShift(BitMask,Int32).right.parameter.Out.0\ <= to_signed(8, 32);
                            \Unum::ExponentSize().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ <= true;
                            \Unum::ExponentSize().0._State\ := \Unum::ExponentSize().0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentSize().0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_RightShift(Lombiq.Unum.BitMask,System.Int32)
                        if (\Unum::ExponentSize().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ = \Unum::ExponentSize().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\) then 
                            \Unum::ExponentSize().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ <= false;
                            \Unum::ExponentSize().0.return.2\ := \Unum::ExponentSize().0.BitMask::op_RightShift(BitMask,Int32).return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,System.UInt32)
                            \Unum::ExponentSize().0.BitMask::op_Addition(BitMask,UInt32).left.parameter.Out.0\ <= \Unum::ExponentSize().0.return.2\;
                            \Unum::ExponentSize().0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\ <= to_unsigned(1, 32);
                            \Unum::ExponentSize().0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ <= true;
                            \Unum::ExponentSize().0._State\ := \Unum::ExponentSize().0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentSize().0._State_6\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,System.UInt32)
                        if (\Unum::ExponentSize().0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ = \Unum::ExponentSize().0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\) then 
                            \Unum::ExponentSize().0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ <= false;
                            \Unum::ExponentSize().0.return.3\ := \Unum::ExponentSize().0.BitMask::op_Addition(BitMask,UInt32).return.0\;
                            -- Starting state machine invocation for the following method: System.UInt32 Lombiq.Unum.BitMask::GetLowest32Bits()
                            \Unum::ExponentSize().0.BitMask::GetLowest32Bits().this.parameter.Out.0\ <= \Unum::ExponentSize().0.return.3\;
                            \Unum::ExponentSize().0.BitMask::GetLowest32Bits()._Started.0\ <= true;
                            \Unum::ExponentSize().0._State\ := \Unum::ExponentSize().0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentSize().0._State_7\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Lombiq.Unum.BitMask::GetLowest32Bits()
                        if (\Unum::ExponentSize().0.BitMask::GetLowest32Bits()._Started.0\ = \Unum::ExponentSize().0.BitMask::GetLowest32Bits()._Finished.0\) then 
                            \Unum::ExponentSize().0.BitMask::GetLowest32Bits()._Started.0\ <= false;
                            \Unum::ExponentSize().0.return.4\ := \Unum::ExponentSize().0.BitMask::GetLowest32Bits().return.0\;
                            \Unum::ExponentSize().0.return\ <= resize(\Unum::ExponentSize().0.return.4\, 8);
                            \Unum::ExponentSize().0._State\ := \Unum::ExponentSize().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Byte Lombiq.Unum.Unum::ExponentSize().0 state machine end


    -- System.UInt16 Lombiq.Unum.Unum::FractionSize().0 state machine start
    \Unum::FractionSize().0._StateMachine\: process (\Clock\) 
        Variable \Unum::FractionSize().0._State\: \Unum::FractionSize().0._States\ := \Unum::FractionSize().0._State_0\;
        Variable \Unum::FractionSize().0.this\: \Lombiq.Unum.Unum\;
        Variable \Unum::FractionSize().0.return.0\: \Lombiq.Unum.BitMask\;
        Variable \Unum::FractionSize().0.return.1\: \Lombiq.Unum.BitMask\;
        Variable \Unum::FractionSize().0.return.2\: \Lombiq.Unum.BitMask\;
        Variable \Unum::FractionSize().0.return.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::FractionSize().0._Finished\ <= false;
                \Unum::FractionSize().0.return\ <= to_unsigned(0, 16);
                \Unum::FractionSize().0.Unum::get_FractionSizeMask()._Started.0\ <= false;
                \Unum::FractionSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ <= false;
                \Unum::FractionSize().0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\ <= to_unsigned(0, 32);
                \Unum::FractionSize().0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ <= false;
                \Unum::FractionSize().0.BitMask::GetLowest32Bits()._Started.0\ <= false;
                \Unum::FractionSize().0._State\ := \Unum::FractionSize().0._State_0\;
                \Unum::FractionSize().0.return.3\ := to_unsigned(0, 32);
            else 
                case \Unum::FractionSize().0._State\ is 
                    when \Unum::FractionSize().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::FractionSize().0._Started\ = true) then 
                            \Unum::FractionSize().0._State\ := \Unum::FractionSize().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionSize().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::FractionSize().0._Started\ = true) then 
                            \Unum::FractionSize().0._Finished\ <= true;
                        else 
                            \Unum::FractionSize().0._Finished\ <= false;
                            \Unum::FractionSize().0._State\ := \Unum::FractionSize().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionSize().0._State_2\ => 
                        \Unum::FractionSize().0.this\ := \Unum::FractionSize().0.this.parameter.In\;
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_FractionSizeMask()
                        \Unum::FractionSize().0.Unum::get_FractionSizeMask().this.parameter.Out.0\ <= \Unum::FractionSize().0.this\;
                        \Unum::FractionSize().0.Unum::get_FractionSizeMask()._Started.0\ <= true;
                        \Unum::FractionSize().0._State\ := \Unum::FractionSize().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionSize().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_FractionSizeMask()
                        if (\Unum::FractionSize().0.Unum::get_FractionSizeMask()._Started.0\ = \Unum::FractionSize().0.Unum::get_FractionSizeMask()._Finished.0\) then 
                            \Unum::FractionSize().0.Unum::get_FractionSizeMask()._Started.0\ <= false;
                            \Unum::FractionSize().0.return.0\ := \Unum::FractionSize().0.Unum::get_FractionSizeMask().return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseAnd(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \Unum::FractionSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask).left.parameter.Out.0\ <= \Unum::FractionSize().0.this\.\UnumBits\;
                            \Unum::FractionSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask).right.parameter.Out.0\ <= \Unum::FractionSize().0.return.0\;
                            \Unum::FractionSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ <= true;
                            \Unum::FractionSize().0._State\ := \Unum::FractionSize().0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionSize().0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseAnd(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\Unum::FractionSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ = \Unum::FractionSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\) then 
                            \Unum::FractionSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ <= false;
                            \Unum::FractionSize().0.return.1\ := \Unum::FractionSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask).return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,System.UInt32)
                            \Unum::FractionSize().0.BitMask::op_Addition(BitMask,UInt32).left.parameter.Out.0\ <= \Unum::FractionSize().0.return.1\;
                            \Unum::FractionSize().0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\ <= to_unsigned(1, 32);
                            \Unum::FractionSize().0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ <= true;
                            \Unum::FractionSize().0._State\ := \Unum::FractionSize().0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionSize().0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,System.UInt32)
                        if (\Unum::FractionSize().0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ = \Unum::FractionSize().0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\) then 
                            \Unum::FractionSize().0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ <= false;
                            \Unum::FractionSize().0.return.2\ := \Unum::FractionSize().0.BitMask::op_Addition(BitMask,UInt32).return.0\;
                            -- Starting state machine invocation for the following method: System.UInt32 Lombiq.Unum.BitMask::GetLowest32Bits()
                            \Unum::FractionSize().0.BitMask::GetLowest32Bits().this.parameter.Out.0\ <= \Unum::FractionSize().0.return.2\;
                            \Unum::FractionSize().0.BitMask::GetLowest32Bits()._Started.0\ <= true;
                            \Unum::FractionSize().0._State\ := \Unum::FractionSize().0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionSize().0._State_6\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Lombiq.Unum.BitMask::GetLowest32Bits()
                        if (\Unum::FractionSize().0.BitMask::GetLowest32Bits()._Started.0\ = \Unum::FractionSize().0.BitMask::GetLowest32Bits()._Finished.0\) then 
                            \Unum::FractionSize().0.BitMask::GetLowest32Bits()._Started.0\ <= false;
                            \Unum::FractionSize().0.return.3\ := \Unum::FractionSize().0.BitMask::GetLowest32Bits().return.0\;
                            \Unum::FractionSize().0.return\ <= resize(\Unum::FractionSize().0.return.3\, 16);
                            \Unum::FractionSize().0._State\ := \Unum::FractionSize().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.UInt16 Lombiq.Unum.Unum::FractionSize().0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionMask().0 state machine start
    \Unum::FractionMask().0._StateMachine\: process (\Clock\) 
        Variable \Unum::FractionMask().0._State\: \Unum::FractionMask().0._States\ := \Unum::FractionMask().0._State_0\;
        Variable \Unum::FractionMask().0.this\: \Lombiq.Unum.Unum\;
        Variable \Unum::FractionMask().0.left\: \Lombiq.Unum.BitMask\;
        Variable \Unum::FractionMask().0.array6d2b985ad94fec35ed2e2f13cc3bf07ded4f1c91959baba527e335c63d6a51ad\: \unsigned32_Array\(0 to 0) := (others => to_unsigned(0, 32));
        Variable \Unum::FractionMask().0.return.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::FractionMask().0.return.1\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::FractionMask().0.return.2\: \Lombiq.Unum.BitMask\;
        Variable \Unum::FractionMask().0.return.3\: \Lombiq.Unum.BitMask\;
        Variable \Unum::FractionMask().0.return.4\: \Lombiq.Unum.BitMask\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::FractionMask().0._Finished\ <= false;
                \Unum::FractionMask().0.Unum::get_Size()._Started.0\ <= false;
                \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 32));
                \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                \Unum::FractionMask().0.Unum::FractionSize()._Started.0\ <= false;
                \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\ <= to_signed(0, 32);
                \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= false;
                \Unum::FractionMask().0.BitMask::op_Subtraction(BitMask,UInt32).right.parameter.Out.0\ <= to_unsigned(0, 32);
                \Unum::FractionMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ <= false;
                \Unum::FractionMask().0._State\ := \Unum::FractionMask().0._State_0\;
                \Unum::FractionMask().0.array6d2b985ad94fec35ed2e2f13cc3bf07ded4f1c91959baba527e335c63d6a51ad\ := (others => to_unsigned(0, 32));
                \Unum::FractionMask().0.return.0\ := to_unsigned(0, 16);
                \Unum::FractionMask().0.return.1\ := to_unsigned(0, 16);
            else 
                case \Unum::FractionMask().0._State\ is 
                    when \Unum::FractionMask().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::FractionMask().0._Started\ = true) then 
                            \Unum::FractionMask().0._State\ := \Unum::FractionMask().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionMask().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::FractionMask().0._Started\ = true) then 
                            \Unum::FractionMask().0._Finished\ <= true;
                        else 
                            \Unum::FractionMask().0._Finished\ <= false;
                            \Unum::FractionMask().0._State\ := \Unum::FractionMask().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionMask().0._State_2\ => 
                        \Unum::FractionMask().0.this\ := \Unum::FractionMask().0.this.parameter.In\;
                        \Unum::FractionMask().0.array6d2b985ad94fec35ed2e2f13cc3bf07ded4f1c91959baba527e335c63d6a51ad\ := (others => to_unsigned(0, 32));
                        \Unum::FractionMask().0.array6d2b985ad94fec35ed2e2f13cc3bf07ded4f1c91959baba527e335c63d6a51ad\(to_integer(to_signed(0, 32))) := to_unsigned(1, 32);
                        -- Initializing record fields to their defaults.
                        \Unum::FractionMask().0.left\.\IsNull\ := false;
                        \Unum::FractionMask().0.left\.\Size\ := to_unsigned(0, 16);
                        \Unum::FractionMask().0.left\.\SegmentCount\ := to_unsigned(0, 16);
                        \Unum::FractionMask().0.left\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::get_Size()
                        \Unum::FractionMask().0.Unum::get_Size().this.parameter.Out.0\ <= \Unum::FractionMask().0.this\;
                        \Unum::FractionMask().0.Unum::get_Size()._Started.0\ <= true;
                        \Unum::FractionMask().0._State\ := \Unum::FractionMask().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionMask().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::get_Size()
                        if (\Unum::FractionMask().0.Unum::get_Size()._Started.0\ = \Unum::FractionMask().0.Unum::get_Size()._Finished.0\) then 
                            \Unum::FractionMask().0.Unum::get_Size()._Started.0\ <= false;
                            \Unum::FractionMask().0.return.0\ := \Unum::FractionMask().0.Unum::get_Size().return.0\;
                            -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                            \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\ <= \Unum::FractionMask().0.left\;
                            \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\(0 to 0) <= \Unum::FractionMask().0.array6d2b985ad94fec35ed2e2f13cc3bf07ded4f1c91959baba527e335c63d6a51ad\;
                            \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= \Unum::FractionMask().0.return.0\;
                            \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= true;
                            \Unum::FractionMask().0._State\ := \Unum::FractionMask().0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionMask().0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        if (\Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\) then 
                            \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                            \Unum::FractionMask().0.left\ := \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\;
                            \Unum::FractionMask().0.array6d2b985ad94fec35ed2e2f13cc3bf07ded4f1c91959baba527e335c63d6a51ad\ := \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\(0 to 0);
                            -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::FractionSize()
                            \Unum::FractionMask().0.Unum::FractionSize()._Started.0\ <= true;
                            \Unum::FractionMask().0._State\ := \Unum::FractionMask().0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionMask().0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::FractionSize()
                        if (\Unum::FractionMask().0.Unum::FractionSize()._Started.0\ = \Unum::FractionMask().0.Unum::FractionSize()._Finished.0\) then 
                            \Unum::FractionMask().0.Unum::FractionSize()._Started.0\ <= false;
                            \Unum::FractionMask().0.return.1\ := \Unum::FractionMask().0.Unum::FractionSize().return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                            \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\ <= \Unum::FractionMask().0.left\;
                            \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\ <= resize(signed(\Unum::FractionMask().0.return.1\), 32);
                            \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= true;
                            \Unum::FractionMask().0._State\ := \Unum::FractionMask().0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionMask().0._State_6\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                        if (\Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ = \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\) then 
                            \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= false;
                            \Unum::FractionMask().0.return.2\ := \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32).return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,System.UInt32)
                            \Unum::FractionMask().0.BitMask::op_Subtraction(BitMask,UInt32).left.parameter.Out.0\ <= \Unum::FractionMask().0.return.2\;
                            \Unum::FractionMask().0.BitMask::op_Subtraction(BitMask,UInt32).right.parameter.Out.0\ <= to_unsigned(1, 32);
                            \Unum::FractionMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ <= true;
                            \Unum::FractionMask().0._State\ := \Unum::FractionMask().0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionMask().0._State_7\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,System.UInt32)
                        if (\Unum::FractionMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ = \Unum::FractionMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\) then 
                            \Unum::FractionMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ <= false;
                            \Unum::FractionMask().0.return.3\ := \Unum::FractionMask().0.BitMask::op_Subtraction(BitMask,UInt32).return.0\;
                            -- The last invocation for the target state machine finished in the previous state, so need to start the next one in the next state.
                            \Unum::FractionMask().0._State\ := \Unum::FractionMask().0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionMask().0._State_8\ => 
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                        \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\ <= \Unum::FractionMask().0.return.3\;
                        \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\ <= to_signed(13, 32);
                        \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= true;
                        \Unum::FractionMask().0._State\ := \Unum::FractionMask().0._State_9\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionMask().0._State_9\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                        if (\Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ = \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\) then 
                            \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= false;
                            \Unum::FractionMask().0.return.4\ := \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32).return.0\;
                            \Unum::FractionMask().0.return\ <= \Unum::FractionMask().0.return.4\;
                            \Unum::FractionMask().0._State\ := \Unum::FractionMask().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionMask().0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentMask().0 state machine start
    \Unum::ExponentMask().0._StateMachine\: process (\Clock\) 
        Variable \Unum::ExponentMask().0._State\: \Unum::ExponentMask().0._States\ := \Unum::ExponentMask().0._State_0\;
        Variable \Unum::ExponentMask().0.this\: \Lombiq.Unum.Unum\;
        Variable \Unum::ExponentMask().0.left\: \Lombiq.Unum.BitMask\;
        Variable \Unum::ExponentMask().0.array1cc7a004cb9772c19b379599c867170bc2486e605fb7c3de94aec89d8c9df458\: \unsigned32_Array\(0 to 0) := (others => to_unsigned(0, 32));
        Variable \Unum::ExponentMask().0.return.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::ExponentMask().0.return.1\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Unum::ExponentMask().0.return.2\: \Lombiq.Unum.BitMask\;
        Variable \Unum::ExponentMask().0.return.3\: \Lombiq.Unum.BitMask\;
        Variable \Unum::ExponentMask().0.return.4\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::ExponentMask().0.binaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::ExponentMask().0.return.5\: \Lombiq.Unum.BitMask\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::ExponentMask().0._Finished\ <= false;
                \Unum::ExponentMask().0.Unum::get_Size()._Started.0\ <= false;
                \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 32));
                \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                \Unum::ExponentMask().0.Unum::ExponentSize()._Started.0\ <= false;
                \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\ <= to_signed(0, 32);
                \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= false;
                \Unum::ExponentMask().0.BitMask::op_Subtraction(BitMask,UInt32).right.parameter.Out.0\ <= to_unsigned(0, 32);
                \Unum::ExponentMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ <= false;
                \Unum::ExponentMask().0.Unum::FractionSize()._Started.0\ <= false;
                \Unum::ExponentMask().0._State\ := \Unum::ExponentMask().0._State_0\;
                \Unum::ExponentMask().0.array1cc7a004cb9772c19b379599c867170bc2486e605fb7c3de94aec89d8c9df458\ := (others => to_unsigned(0, 32));
                \Unum::ExponentMask().0.return.0\ := to_unsigned(0, 16);
                \Unum::ExponentMask().0.return.1\ := to_unsigned(0, 8);
                \Unum::ExponentMask().0.return.4\ := to_unsigned(0, 16);
                \Unum::ExponentMask().0.binaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \Unum::ExponentMask().0._State\ is 
                    when \Unum::ExponentMask().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::ExponentMask().0._Started\ = true) then 
                            \Unum::ExponentMask().0._State\ := \Unum::ExponentMask().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentMask().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::ExponentMask().0._Started\ = true) then 
                            \Unum::ExponentMask().0._Finished\ <= true;
                        else 
                            \Unum::ExponentMask().0._Finished\ <= false;
                            \Unum::ExponentMask().0._State\ := \Unum::ExponentMask().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentMask().0._State_2\ => 
                        \Unum::ExponentMask().0.this\ := \Unum::ExponentMask().0.this.parameter.In\;
                        \Unum::ExponentMask().0.array1cc7a004cb9772c19b379599c867170bc2486e605fb7c3de94aec89d8c9df458\ := (others => to_unsigned(0, 32));
                        \Unum::ExponentMask().0.array1cc7a004cb9772c19b379599c867170bc2486e605fb7c3de94aec89d8c9df458\(to_integer(to_signed(0, 32))) := to_unsigned(1, 32);
                        -- Initializing record fields to their defaults.
                        \Unum::ExponentMask().0.left\.\IsNull\ := false;
                        \Unum::ExponentMask().0.left\.\Size\ := to_unsigned(0, 16);
                        \Unum::ExponentMask().0.left\.\SegmentCount\ := to_unsigned(0, 16);
                        \Unum::ExponentMask().0.left\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::get_Size()
                        \Unum::ExponentMask().0.Unum::get_Size().this.parameter.Out.0\ <= \Unum::ExponentMask().0.this\;
                        \Unum::ExponentMask().0.Unum::get_Size()._Started.0\ <= true;
                        \Unum::ExponentMask().0._State\ := \Unum::ExponentMask().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentMask().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::get_Size()
                        if (\Unum::ExponentMask().0.Unum::get_Size()._Started.0\ = \Unum::ExponentMask().0.Unum::get_Size()._Finished.0\) then 
                            \Unum::ExponentMask().0.Unum::get_Size()._Started.0\ <= false;
                            \Unum::ExponentMask().0.return.0\ := \Unum::ExponentMask().0.Unum::get_Size().return.0\;
                            -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                            \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\ <= \Unum::ExponentMask().0.left\;
                            \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\(0 to 0) <= \Unum::ExponentMask().0.array1cc7a004cb9772c19b379599c867170bc2486e605fb7c3de94aec89d8c9df458\;
                            \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= \Unum::ExponentMask().0.return.0\;
                            \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= true;
                            \Unum::ExponentMask().0._State\ := \Unum::ExponentMask().0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentMask().0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        if (\Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\) then 
                            \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                            \Unum::ExponentMask().0.left\ := \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\;
                            \Unum::ExponentMask().0.array1cc7a004cb9772c19b379599c867170bc2486e605fb7c3de94aec89d8c9df458\ := \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\(0 to 0);
                            -- Starting state machine invocation for the following method: System.Byte Lombiq.Unum.Unum::ExponentSize()
                            \Unum::ExponentMask().0.Unum::ExponentSize()._Started.0\ <= true;
                            \Unum::ExponentMask().0._State\ := \Unum::ExponentMask().0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentMask().0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Byte Lombiq.Unum.Unum::ExponentSize()
                        if (\Unum::ExponentMask().0.Unum::ExponentSize()._Started.0\ = \Unum::ExponentMask().0.Unum::ExponentSize()._Finished.0\) then 
                            \Unum::ExponentMask().0.Unum::ExponentSize()._Started.0\ <= false;
                            \Unum::ExponentMask().0.return.1\ := \Unum::ExponentMask().0.Unum::ExponentSize().return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                            \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\ <= \Unum::ExponentMask().0.left\;
                            \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\ <= resize(signed(\Unum::ExponentMask().0.return.1\), 32);
                            \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= true;
                            \Unum::ExponentMask().0._State\ := \Unum::ExponentMask().0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentMask().0._State_6\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                        if (\Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ = \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\) then 
                            \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= false;
                            \Unum::ExponentMask().0.return.2\ := \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32).return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,System.UInt32)
                            \Unum::ExponentMask().0.BitMask::op_Subtraction(BitMask,UInt32).left.parameter.Out.0\ <= \Unum::ExponentMask().0.return.2\;
                            \Unum::ExponentMask().0.BitMask::op_Subtraction(BitMask,UInt32).right.parameter.Out.0\ <= to_unsigned(1, 32);
                            \Unum::ExponentMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ <= true;
                            \Unum::ExponentMask().0._State\ := \Unum::ExponentMask().0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentMask().0._State_7\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,System.UInt32)
                        if (\Unum::ExponentMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ = \Unum::ExponentMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\) then 
                            \Unum::ExponentMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ <= false;
                            \Unum::ExponentMask().0.return.3\ := \Unum::ExponentMask().0.BitMask::op_Subtraction(BitMask,UInt32).return.0\;
                            -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::FractionSize()
                            \Unum::ExponentMask().0.Unum::FractionSize()._Started.0\ <= true;
                            \Unum::ExponentMask().0._State\ := \Unum::ExponentMask().0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentMask().0._State_8\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::FractionSize()
                        if (\Unum::ExponentMask().0.Unum::FractionSize()._Started.0\ = \Unum::ExponentMask().0.Unum::FractionSize()._Finished.0\) then 
                            \Unum::ExponentMask().0.Unum::FractionSize()._Started.0\ <= false;
                            \Unum::ExponentMask().0.return.4\ := \Unum::ExponentMask().0.Unum::FractionSize().return.0\;
                            \Unum::ExponentMask().0.binaryOperationResult.0\ := resize(signed(\Unum::ExponentMask().0.return.4\ + to_unsigned(13, 16)), 32);
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                            \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\ <= \Unum::ExponentMask().0.return.3\;
                            \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\ <= (\Unum::ExponentMask().0.binaryOperationResult.0\);
                            \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= true;
                            \Unum::ExponentMask().0._State\ := \Unum::ExponentMask().0._State_9\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::ExponentMask().0._State_9\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                        if (\Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ = \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\) then 
                            \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= false;
                            \Unum::ExponentMask().0.return.5\ := \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32).return.0\;
                            \Unum::ExponentMask().0.return\ <= \Unum::ExponentMask().0.return.5\;
                            \Unum::ExponentMask().0._State\ := \Unum::ExponentMask().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentMask().0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::Exponent().0 state machine start
    \Unum::Exponent().0._StateMachine\: process (\Clock\) 
        Variable \Unum::Exponent().0._State\: \Unum::Exponent().0._States\ := \Unum::Exponent().0._State_0\;
        Variable \Unum::Exponent().0.this\: \Lombiq.Unum.Unum\;
        Variable \Unum::Exponent().0.return.0\: \Lombiq.Unum.BitMask\;
        Variable \Unum::Exponent().0.return.1\: \Lombiq.Unum.BitMask\;
        Variable \Unum::Exponent().0.return.2\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::Exponent().0.binaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::Exponent().0.return.3\: \Lombiq.Unum.BitMask\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::Exponent().0._Finished\ <= false;
                \Unum::Exponent().0.Unum::ExponentMask()._Started.0\ <= false;
                \Unum::Exponent().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ <= false;
                \Unum::Exponent().0.Unum::FractionSize()._Started.0\ <= false;
                \Unum::Exponent().0.BitMask::op_RightShift(BitMask,Int32).right.parameter.Out.0\ <= to_signed(0, 32);
                \Unum::Exponent().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ <= false;
                \Unum::Exponent().0._State\ := \Unum::Exponent().0._State_0\;
                \Unum::Exponent().0.return.2\ := to_unsigned(0, 16);
                \Unum::Exponent().0.binaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \Unum::Exponent().0._State\ is 
                    when \Unum::Exponent().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::Exponent().0._Started\ = true) then 
                            \Unum::Exponent().0._State\ := \Unum::Exponent().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::Exponent().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::Exponent().0._Started\ = true) then 
                            \Unum::Exponent().0._Finished\ <= true;
                        else 
                            \Unum::Exponent().0._Finished\ <= false;
                            \Unum::Exponent().0._State\ := \Unum::Exponent().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::Exponent().0._State_2\ => 
                        \Unum::Exponent().0.this\ := \Unum::Exponent().0.this.parameter.In\;
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentMask()
                        \Unum::Exponent().0.Unum::ExponentMask()._Started.0\ <= true;
                        \Unum::Exponent().0._State\ := \Unum::Exponent().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::Exponent().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentMask()
                        if (\Unum::Exponent().0.Unum::ExponentMask()._Started.0\ = \Unum::Exponent().0.Unum::ExponentMask()._Finished.0\) then 
                            \Unum::Exponent().0.Unum::ExponentMask()._Started.0\ <= false;
                            \Unum::Exponent().0.return.0\ := \Unum::Exponent().0.Unum::ExponentMask().return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseAnd(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \Unum::Exponent().0.BitMask::op_BitwiseAnd(BitMask,BitMask).left.parameter.Out.0\ <= \Unum::Exponent().0.return.0\;
                            \Unum::Exponent().0.BitMask::op_BitwiseAnd(BitMask,BitMask).right.parameter.Out.0\ <= \Unum::Exponent().0.this\.\UnumBits\;
                            \Unum::Exponent().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ <= true;
                            \Unum::Exponent().0._State\ := \Unum::Exponent().0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::Exponent().0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseAnd(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\Unum::Exponent().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ = \Unum::Exponent().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\) then 
                            \Unum::Exponent().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ <= false;
                            \Unum::Exponent().0.return.1\ := \Unum::Exponent().0.BitMask::op_BitwiseAnd(BitMask,BitMask).return.0\;
                            -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::FractionSize()
                            \Unum::Exponent().0.Unum::FractionSize()._Started.0\ <= true;
                            \Unum::Exponent().0._State\ := \Unum::Exponent().0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::Exponent().0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::FractionSize()
                        if (\Unum::Exponent().0.Unum::FractionSize()._Started.0\ = \Unum::Exponent().0.Unum::FractionSize()._Finished.0\) then 
                            \Unum::Exponent().0.Unum::FractionSize()._Started.0\ <= false;
                            \Unum::Exponent().0.return.2\ := \Unum::Exponent().0.Unum::FractionSize().return.0\;
                            \Unum::Exponent().0.binaryOperationResult.0\ := resize(signed(to_unsigned(13, 16) + \Unum::Exponent().0.return.2\), 32);
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_RightShift(Lombiq.Unum.BitMask,System.Int32)
                            \Unum::Exponent().0.BitMask::op_RightShift(BitMask,Int32).left.parameter.Out.0\ <= \Unum::Exponent().0.return.1\;
                            \Unum::Exponent().0.BitMask::op_RightShift(BitMask,Int32).right.parameter.Out.0\ <= (\Unum::Exponent().0.binaryOperationResult.0\);
                            \Unum::Exponent().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ <= true;
                            \Unum::Exponent().0._State\ := \Unum::Exponent().0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::Exponent().0._State_6\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_RightShift(Lombiq.Unum.BitMask,System.Int32)
                        if (\Unum::Exponent().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ = \Unum::Exponent().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\) then 
                            \Unum::Exponent().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ <= false;
                            \Unum::Exponent().0.return.3\ := \Unum::Exponent().0.BitMask::op_RightShift(BitMask,Int32).return.0\;
                            \Unum::Exponent().0.return\ <= \Unum::Exponent().0.return.3\;
                            \Unum::Exponent().0._State\ := \Unum::Exponent().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::Exponent().0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::Fraction().0 state machine start
    \Unum::Fraction().0._StateMachine\: process (\Clock\) 
        Variable \Unum::Fraction().0._State\: \Unum::Fraction().0._States\ := \Unum::Fraction().0._State_0\;
        Variable \Unum::Fraction().0.this\: \Lombiq.Unum.Unum\;
        Variable \Unum::Fraction().0.return.0\: \Lombiq.Unum.BitMask\;
        Variable \Unum::Fraction().0.return.1\: \Lombiq.Unum.BitMask\;
        Variable \Unum::Fraction().0.return.2\: \Lombiq.Unum.BitMask\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::Fraction().0._Finished\ <= false;
                \Unum::Fraction().0.Unum::FractionMask()._Started.0\ <= false;
                \Unum::Fraction().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ <= false;
                \Unum::Fraction().0.BitMask::op_RightShift(BitMask,Int32).right.parameter.Out.0\ <= to_signed(0, 32);
                \Unum::Fraction().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ <= false;
                \Unum::Fraction().0._State\ := \Unum::Fraction().0._State_0\;
            else 
                case \Unum::Fraction().0._State\ is 
                    when \Unum::Fraction().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::Fraction().0._Started\ = true) then 
                            \Unum::Fraction().0._State\ := \Unum::Fraction().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::Fraction().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::Fraction().0._Started\ = true) then 
                            \Unum::Fraction().0._Finished\ <= true;
                        else 
                            \Unum::Fraction().0._Finished\ <= false;
                            \Unum::Fraction().0._State\ := \Unum::Fraction().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::Fraction().0._State_2\ => 
                        \Unum::Fraction().0.this\ := \Unum::Fraction().0.this.parameter.In\;
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionMask()
                        \Unum::Fraction().0.Unum::FractionMask()._Started.0\ <= true;
                        \Unum::Fraction().0._State\ := \Unum::Fraction().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::Fraction().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionMask()
                        if (\Unum::Fraction().0.Unum::FractionMask()._Started.0\ = \Unum::Fraction().0.Unum::FractionMask()._Finished.0\) then 
                            \Unum::Fraction().0.Unum::FractionMask()._Started.0\ <= false;
                            \Unum::Fraction().0.return.0\ := \Unum::Fraction().0.Unum::FractionMask().return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseAnd(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \Unum::Fraction().0.BitMask::op_BitwiseAnd(BitMask,BitMask).left.parameter.Out.0\ <= \Unum::Fraction().0.return.0\;
                            \Unum::Fraction().0.BitMask::op_BitwiseAnd(BitMask,BitMask).right.parameter.Out.0\ <= \Unum::Fraction().0.this\.\UnumBits\;
                            \Unum::Fraction().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ <= true;
                            \Unum::Fraction().0._State\ := \Unum::Fraction().0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::Fraction().0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseAnd(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\Unum::Fraction().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ = \Unum::Fraction().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\) then 
                            \Unum::Fraction().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ <= false;
                            \Unum::Fraction().0.return.1\ := \Unum::Fraction().0.BitMask::op_BitwiseAnd(BitMask,BitMask).return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_RightShift(Lombiq.Unum.BitMask,System.Int32)
                            \Unum::Fraction().0.BitMask::op_RightShift(BitMask,Int32).left.parameter.Out.0\ <= \Unum::Fraction().0.return.1\;
                            \Unum::Fraction().0.BitMask::op_RightShift(BitMask,Int32).right.parameter.Out.0\ <= to_signed(13, 32);
                            \Unum::Fraction().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ <= true;
                            \Unum::Fraction().0._State\ := \Unum::Fraction().0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::Fraction().0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_RightShift(Lombiq.Unum.BitMask,System.Int32)
                        if (\Unum::Fraction().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ = \Unum::Fraction().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\) then 
                            \Unum::Fraction().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ <= false;
                            \Unum::Fraction().0.return.2\ := \Unum::Fraction().0.BitMask::op_RightShift(BitMask,Int32).return.0\;
                            \Unum::Fraction().0.return\ <= \Unum::Fraction().0.return.2\;
                            \Unum::Fraction().0._State\ := \Unum::Fraction().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::Fraction().0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit().0 state machine start
    \Unum::FractionWithHiddenBit().0._StateMachine\: process (\Clock\) 
        Variable \Unum::FractionWithHiddenBit().0._State\: \Unum::FractionWithHiddenBit().0._States\ := \Unum::FractionWithHiddenBit().0._State_0\;
        Variable \Unum::FractionWithHiddenBit().0.this\: \Lombiq.Unum.Unum\;
        Variable \Unum::FractionWithHiddenBit().0.conditionald0fe2758c76631203a5f7ea7a5ba0e2f98df065961f41fa3c746fb0d250f2d75\: \Lombiq.Unum.BitMask\;
        Variable \Unum::FractionWithHiddenBit().0.return.0\: boolean := false;
        Variable \Unum::FractionWithHiddenBit().0.return.1\: \Lombiq.Unum.BitMask\;
        Variable \Unum::FractionWithHiddenBit().0.return.2\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::FractionWithHiddenBit().0.return.3\: \Lombiq.Unum.BitMask\;
        Variable \Unum::FractionWithHiddenBit().0.return.4\: \Lombiq.Unum.BitMask\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::FractionWithHiddenBit().0._Finished\ <= false;
                \Unum::FractionWithHiddenBit().0.Unum::HiddenBitIsOne()._Started.0\ <= false;
                \Unum::FractionWithHiddenBit().0.Unum::Fraction()._Started.0\ <= false;
                \Unum::FractionWithHiddenBit().0.Unum::FractionSize()._Started.0\ <= false;
                \Unum::FractionWithHiddenBit().0.BitMask::SetOne(UInt16).index.parameter.Out.0\ <= to_unsigned(0, 16);
                \Unum::FractionWithHiddenBit().0.BitMask::SetOne(UInt16)._Started.0\ <= false;
                \Unum::FractionWithHiddenBit().0._State\ := \Unum::FractionWithHiddenBit().0._State_0\;
                \Unum::FractionWithHiddenBit().0.return.0\ := false;
                \Unum::FractionWithHiddenBit().0.return.2\ := to_unsigned(0, 16);
            else 
                case \Unum::FractionWithHiddenBit().0._State\ is 
                    when \Unum::FractionWithHiddenBit().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::FractionWithHiddenBit().0._Started\ = true) then 
                            \Unum::FractionWithHiddenBit().0._State\ := \Unum::FractionWithHiddenBit().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionWithHiddenBit().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::FractionWithHiddenBit().0._Started\ = true) then 
                            \Unum::FractionWithHiddenBit().0._Finished\ <= true;
                        else 
                            \Unum::FractionWithHiddenBit().0._Finished\ <= false;
                            \Unum::FractionWithHiddenBit().0._State\ := \Unum::FractionWithHiddenBit().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionWithHiddenBit().0._State_2\ => 
                        \Unum::FractionWithHiddenBit().0.this\ := \Unum::FractionWithHiddenBit().0.this.parameter.In\;
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::HiddenBitIsOne()
                        \Unum::FractionWithHiddenBit().0.Unum::HiddenBitIsOne().this.parameter.Out.0\ <= \Unum::FractionWithHiddenBit().0.this\;
                        \Unum::FractionWithHiddenBit().0.Unum::HiddenBitIsOne()._Started.0\ <= true;
                        \Unum::FractionWithHiddenBit().0._State\ := \Unum::FractionWithHiddenBit().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionWithHiddenBit().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::HiddenBitIsOne()
                        if (\Unum::FractionWithHiddenBit().0.Unum::HiddenBitIsOne()._Started.0\ = \Unum::FractionWithHiddenBit().0.Unum::HiddenBitIsOne()._Finished.0\) then 
                            \Unum::FractionWithHiddenBit().0.Unum::HiddenBitIsOne()._Started.0\ <= false;
                            \Unum::FractionWithHiddenBit().0.return.0\ := \Unum::FractionWithHiddenBit().0.Unum::HiddenBitIsOne().return.0\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::FractionWithHiddenBit().0._State_5\ and ends in state \Unum::FractionWithHiddenBit().0._State_8\.
                            --     * The false branch starts in state \Unum::FractionWithHiddenBit().0._State_9\ and ends in state \Unum::FractionWithHiddenBit().0._State_10\.
                            --     * Execution after either branch will continue in the following state: \Unum::FractionWithHiddenBit().0._State_4\.

                            if (\Unum::FractionWithHiddenBit().0.return.0\) then 
                                \Unum::FractionWithHiddenBit().0._State\ := \Unum::FractionWithHiddenBit().0._State_5\;
                            else 
                                \Unum::FractionWithHiddenBit().0._State\ := \Unum::FractionWithHiddenBit().0._State_9\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionWithHiddenBit().0._State_4\ => 
                        -- State after the if-else which was started in state \Unum::FractionWithHiddenBit().0._State_3\.
                        \Unum::FractionWithHiddenBit().0.return\ <= \Unum::FractionWithHiddenBit().0.conditionald0fe2758c76631203a5f7ea7a5ba0e2f98df065961f41fa3c746fb0d250f2d75\;
                        \Unum::FractionWithHiddenBit().0._State\ := \Unum::FractionWithHiddenBit().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionWithHiddenBit().0._State_5\ => 
                        -- True branch of the if-else started in state \Unum::FractionWithHiddenBit().0._State_3\.
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::Fraction()
                        \Unum::FractionWithHiddenBit().0.Unum::Fraction()._Started.0\ <= true;
                        \Unum::FractionWithHiddenBit().0._State\ := \Unum::FractionWithHiddenBit().0._State_6\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionWithHiddenBit().0._State_6\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::Fraction()
                        if (\Unum::FractionWithHiddenBit().0.Unum::Fraction()._Started.0\ = \Unum::FractionWithHiddenBit().0.Unum::Fraction()._Finished.0\) then 
                            \Unum::FractionWithHiddenBit().0.Unum::Fraction()._Started.0\ <= false;
                            \Unum::FractionWithHiddenBit().0.return.1\ := \Unum::FractionWithHiddenBit().0.Unum::Fraction().return.0\;
                            -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::FractionSize()
                            \Unum::FractionWithHiddenBit().0.Unum::FractionSize()._Started.0\ <= true;
                            \Unum::FractionWithHiddenBit().0._State\ := \Unum::FractionWithHiddenBit().0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionWithHiddenBit().0._State_7\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::FractionSize()
                        if (\Unum::FractionWithHiddenBit().0.Unum::FractionSize()._Started.0\ = \Unum::FractionWithHiddenBit().0.Unum::FractionSize()._Finished.0\) then 
                            \Unum::FractionWithHiddenBit().0.Unum::FractionSize()._Started.0\ <= false;
                            \Unum::FractionWithHiddenBit().0.return.2\ := \Unum::FractionWithHiddenBit().0.Unum::FractionSize().return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetOne(System.UInt16)
                            \Unum::FractionWithHiddenBit().0.BitMask::SetOne(UInt16).this.parameter.Out.0\ <= \Unum::FractionWithHiddenBit().0.return.1\;
                            \Unum::FractionWithHiddenBit().0.BitMask::SetOne(UInt16).index.parameter.Out.0\ <= \Unum::FractionWithHiddenBit().0.return.2\;
                            \Unum::FractionWithHiddenBit().0.BitMask::SetOne(UInt16)._Started.0\ <= true;
                            \Unum::FractionWithHiddenBit().0._State\ := \Unum::FractionWithHiddenBit().0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionWithHiddenBit().0._State_8\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetOne(System.UInt16)
                        if (\Unum::FractionWithHiddenBit().0.BitMask::SetOne(UInt16)._Started.0\ = \Unum::FractionWithHiddenBit().0.BitMask::SetOne(UInt16)._Finished.0\) then 
                            \Unum::FractionWithHiddenBit().0.BitMask::SetOne(UInt16)._Started.0\ <= false;
                            \Unum::FractionWithHiddenBit().0.return.3\ := \Unum::FractionWithHiddenBit().0.BitMask::SetOne(UInt16).return.0\;
                            \Unum::FractionWithHiddenBit().0.conditionald0fe2758c76631203a5f7ea7a5ba0e2f98df065961f41fa3c746fb0d250f2d75\ := \Unum::FractionWithHiddenBit().0.return.3\;
                            -- Going to the state after the if-else which was started in state \Unum::FractionWithHiddenBit().0._State_3\.
                            if (\Unum::FractionWithHiddenBit().0._State\ = \Unum::FractionWithHiddenBit().0._State_8\) then 
                                \Unum::FractionWithHiddenBit().0._State\ := \Unum::FractionWithHiddenBit().0._State_4\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionWithHiddenBit().0._State_9\ => 
                        -- False branch of the if-else started in state \Unum::FractionWithHiddenBit().0._State_3\.
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::Fraction()
                        \Unum::FractionWithHiddenBit().0.Unum::Fraction()._Started.0\ <= true;
                        \Unum::FractionWithHiddenBit().0._State\ := \Unum::FractionWithHiddenBit().0._State_10\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::FractionWithHiddenBit().0._State_10\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::Fraction()
                        if (\Unum::FractionWithHiddenBit().0.Unum::Fraction()._Started.0\ = \Unum::FractionWithHiddenBit().0.Unum::Fraction()._Finished.0\) then 
                            \Unum::FractionWithHiddenBit().0.Unum::Fraction()._Started.0\ <= false;
                            \Unum::FractionWithHiddenBit().0.return.4\ := \Unum::FractionWithHiddenBit().0.Unum::Fraction().return.0\;
                            \Unum::FractionWithHiddenBit().0.conditionald0fe2758c76631203a5f7ea7a5ba0e2f98df065961f41fa3c746fb0d250f2d75\ := \Unum::FractionWithHiddenBit().0.return.4\;
                            -- Going to the state after the if-else which was started in state \Unum::FractionWithHiddenBit().0._State_3\.
                            if (\Unum::FractionWithHiddenBit().0._State\ = \Unum::FractionWithHiddenBit().0._State_10\) then 
                                \Unum::FractionWithHiddenBit().0._State\ := \Unum::FractionWithHiddenBit().0._State_4\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit().0 state machine end


    -- System.Int32 Lombiq.Unum.Unum::Bias().0 state machine start
    \Unum::Bias().0._StateMachine\: process (\Clock\) 
        Variable \Unum::Bias().0._State\: \Unum::Bias().0._States\ := \Unum::Bias().0._State_0\;
        Variable \Unum::Bias().0.this\: \Lombiq.Unum.Unum\;
        Variable \Unum::Bias().0.return.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Unum::Bias().0.binaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::Bias().0.binaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::Bias().0.binaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::Bias().0._Finished\ <= false;
                \Unum::Bias().0.return\ <= to_signed(0, 32);
                \Unum::Bias().0.Unum::ExponentSize()._Started.0\ <= false;
                \Unum::Bias().0._State\ := \Unum::Bias().0._State_0\;
                \Unum::Bias().0.return.0\ := to_unsigned(0, 8);
                \Unum::Bias().0.binaryOperationResult.0\ := to_signed(0, 32);
                \Unum::Bias().0.binaryOperationResult.1\ := to_signed(0, 32);
                \Unum::Bias().0.binaryOperationResult.2\ := to_signed(0, 32);
            else 
                case \Unum::Bias().0._State\ is 
                    when \Unum::Bias().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::Bias().0._Started\ = true) then 
                            \Unum::Bias().0._State\ := \Unum::Bias().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::Bias().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::Bias().0._Started\ = true) then 
                            \Unum::Bias().0._Finished\ <= true;
                        else 
                            \Unum::Bias().0._Finished\ <= false;
                            \Unum::Bias().0._State\ := \Unum::Bias().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::Bias().0._State_2\ => 
                        \Unum::Bias().0.this\ := \Unum::Bias().0.this.parameter.In\;
                        -- Starting state machine invocation for the following method: System.Byte Lombiq.Unum.Unum::ExponentSize()
                        \Unum::Bias().0.Unum::ExponentSize()._Started.0\ <= true;
                        \Unum::Bias().0._State\ := \Unum::Bias().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::Bias().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Byte Lombiq.Unum.Unum::ExponentSize()
                        if (\Unum::Bias().0.Unum::ExponentSize()._Started.0\ = \Unum::Bias().0.Unum::ExponentSize()._Finished.0\) then 
                            \Unum::Bias().0.Unum::ExponentSize()._Started.0\ <= false;
                            \Unum::Bias().0.return.0\ := \Unum::Bias().0.Unum::ExponentSize().return.0\;
                            \Unum::Bias().0.binaryOperationResult.0\ := resize(signed(\Unum::Bias().0.return.0\ - to_unsigned(1, 8)), 32);
                            \Unum::Bias().0.binaryOperationResult.1\ := resize(shift_left(to_signed(1, 32), to_integer((\Unum::Bias().0.binaryOperationResult.0\))), 32);
                            \Unum::Bias().0.binaryOperationResult.2\ := \Unum::Bias().0.binaryOperationResult.1\ - to_signed(1, 32);
                            \Unum::Bias().0.return\ <= \Unum::Bias().0.binaryOperationResult.2\;
                            \Unum::Bias().0._State\ := \Unum::Bias().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                end case;
            end if;
        end if;
    end process;
    -- System.Int32 Lombiq.Unum.Unum::Bias().0 state machine end


    -- System.Boolean Lombiq.Unum.Unum::HiddenBitIsOne().0 state machine start
    \Unum::HiddenBitIsOne().0._StateMachine\: process (\Clock\) 
        Variable \Unum::HiddenBitIsOne().0._State\: \Unum::HiddenBitIsOne().0._States\ := \Unum::HiddenBitIsOne().0._State_0\;
        Variable \Unum::HiddenBitIsOne().0.this\: \Lombiq.Unum.Unum\;
        Variable \Unum::HiddenBitIsOne().0.return.0\: \Lombiq.Unum.BitMask\;
        Variable \Unum::HiddenBitIsOne().0.return.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Unum::HiddenBitIsOne().0.binaryOperationResult.0\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::HiddenBitIsOne().0._Finished\ <= false;
                \Unum::HiddenBitIsOne().0.return\ <= false;
                \Unum::HiddenBitIsOne().0.Unum::Exponent()._Started.0\ <= false;
                \Unum::HiddenBitIsOne().0.BitMask::GetLowest32Bits()._Started.0\ <= false;
                \Unum::HiddenBitIsOne().0._State\ := \Unum::HiddenBitIsOne().0._State_0\;
                \Unum::HiddenBitIsOne().0.return.1\ := to_unsigned(0, 32);
                \Unum::HiddenBitIsOne().0.binaryOperationResult.0\ := false;
            else 
                case \Unum::HiddenBitIsOne().0._State\ is 
                    when \Unum::HiddenBitIsOne().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::HiddenBitIsOne().0._Started\ = true) then 
                            \Unum::HiddenBitIsOne().0._State\ := \Unum::HiddenBitIsOne().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::HiddenBitIsOne().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::HiddenBitIsOne().0._Started\ = true) then 
                            \Unum::HiddenBitIsOne().0._Finished\ <= true;
                        else 
                            \Unum::HiddenBitIsOne().0._Finished\ <= false;
                            \Unum::HiddenBitIsOne().0._State\ := \Unum::HiddenBitIsOne().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::HiddenBitIsOne().0._State_2\ => 
                        \Unum::HiddenBitIsOne().0.this\ := \Unum::HiddenBitIsOne().0.this.parameter.In\;
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::Exponent()
                        \Unum::HiddenBitIsOne().0.Unum::Exponent()._Started.0\ <= true;
                        \Unum::HiddenBitIsOne().0._State\ := \Unum::HiddenBitIsOne().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::HiddenBitIsOne().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::Exponent()
                        if (\Unum::HiddenBitIsOne().0.Unum::Exponent()._Started.0\ = \Unum::HiddenBitIsOne().0.Unum::Exponent()._Finished.0\) then 
                            \Unum::HiddenBitIsOne().0.Unum::Exponent()._Started.0\ <= false;
                            \Unum::HiddenBitIsOne().0.return.0\ := \Unum::HiddenBitIsOne().0.Unum::Exponent().return.0\;
                            -- Starting state machine invocation for the following method: System.UInt32 Lombiq.Unum.BitMask::GetLowest32Bits()
                            \Unum::HiddenBitIsOne().0.BitMask::GetLowest32Bits().this.parameter.Out.0\ <= \Unum::HiddenBitIsOne().0.return.0\;
                            \Unum::HiddenBitIsOne().0.BitMask::GetLowest32Bits()._Started.0\ <= true;
                            \Unum::HiddenBitIsOne().0._State\ := \Unum::HiddenBitIsOne().0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::HiddenBitIsOne().0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Lombiq.Unum.BitMask::GetLowest32Bits()
                        if (\Unum::HiddenBitIsOne().0.BitMask::GetLowest32Bits()._Started.0\ = \Unum::HiddenBitIsOne().0.BitMask::GetLowest32Bits()._Finished.0\) then 
                            \Unum::HiddenBitIsOne().0.BitMask::GetLowest32Bits()._Started.0\ <= false;
                            \Unum::HiddenBitIsOne().0.return.1\ := \Unum::HiddenBitIsOne().0.BitMask::GetLowest32Bits().return.0\;
                            \Unum::HiddenBitIsOne().0.binaryOperationResult.0\ := \Unum::HiddenBitIsOne().0.return.1\ > to_unsigned(0, 32);
                            \Unum::HiddenBitIsOne().0.return\ <= \Unum::HiddenBitIsOne().0.binaryOperationResult.0\;
                            \Unum::HiddenBitIsOne().0._State\ := \Unum::HiddenBitIsOne().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Lombiq.Unum.Unum::HiddenBitIsOne().0 state machine end


    -- System.Int32 Lombiq.Unum.Unum::ExponentValueWithBias().0 state machine start
    \Unum::ExponentValueWithBias().0._StateMachine\: process (\Clock\) 
        Variable \Unum::ExponentValueWithBias().0._State\: \Unum::ExponentValueWithBias().0._States\ := \Unum::ExponentValueWithBias().0._State_0\;
        Variable \Unum::ExponentValueWithBias().0.this\: \Lombiq.Unum.Unum\;
        Variable \Unum::ExponentValueWithBias().0.conditional45e7bd3495aef0adb29743d60986bee4963f49e22dbfea77daec45939a162bd1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Unum::ExponentValueWithBias().0.return.0\: boolean := false;
        Variable \Unum::ExponentValueWithBias().0.return.1\: \Lombiq.Unum.BitMask\;
        Variable \Unum::ExponentValueWithBias().0.return.2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Unum::ExponentValueWithBias().0.return.3\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::ExponentValueWithBias().0.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Unum::ExponentValueWithBias().0.binaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::ExponentValueWithBias().0._Finished\ <= false;
                \Unum::ExponentValueWithBias().0.return\ <= to_signed(0, 32);
                \Unum::ExponentValueWithBias().0.Unum::HiddenBitIsOne()._Started.0\ <= false;
                \Unum::ExponentValueWithBias().0.Unum::Exponent()._Started.0\ <= false;
                \Unum::ExponentValueWithBias().0.BitMask::GetLowest32Bits()._Started.0\ <= false;
                \Unum::ExponentValueWithBias().0.Unum::Bias()._Started.0\ <= false;
                \Unum::ExponentValueWithBias().0._State\ := \Unum::ExponentValueWithBias().0._State_0\;
                \Unum::ExponentValueWithBias().0.conditional45e7bd3495aef0adb29743d60986bee4963f49e22dbfea77daec45939a162bd1\ := to_unsigned(0, 32);
                \Unum::ExponentValueWithBias().0.return.0\ := false;
                \Unum::ExponentValueWithBias().0.return.2\ := to_unsigned(0, 32);
                \Unum::ExponentValueWithBias().0.return.3\ := to_signed(0, 32);
                \Unum::ExponentValueWithBias().0.binaryOperationResult.0\ := to_unsigned(0, 32);
                \Unum::ExponentValueWithBias().0.binaryOperationResult.1\ := to_signed(0, 32);
            else 
                case \Unum::ExponentValueWithBias().0._State\ is 
                    when \Unum::ExponentValueWithBias().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::ExponentValueWithBias().0._Started\ = true) then 
                            \Unum::ExponentValueWithBias().0._State\ := \Unum::ExponentValueWithBias().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentValueWithBias().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::ExponentValueWithBias().0._Started\ = true) then 
                            \Unum::ExponentValueWithBias().0._Finished\ <= true;
                        else 
                            \Unum::ExponentValueWithBias().0._Finished\ <= false;
                            \Unum::ExponentValueWithBias().0._State\ := \Unum::ExponentValueWithBias().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentValueWithBias().0._State_2\ => 
                        \Unum::ExponentValueWithBias().0.this\ := \Unum::ExponentValueWithBias().0.this.parameter.In\;
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::HiddenBitIsOne()
                        \Unum::ExponentValueWithBias().0.Unum::HiddenBitIsOne()._Started.0\ <= true;
                        \Unum::ExponentValueWithBias().0._State\ := \Unum::ExponentValueWithBias().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentValueWithBias().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::HiddenBitIsOne()
                        if (\Unum::ExponentValueWithBias().0.Unum::HiddenBitIsOne()._Started.0\ = \Unum::ExponentValueWithBias().0.Unum::HiddenBitIsOne()._Finished.0\) then 
                            \Unum::ExponentValueWithBias().0.Unum::HiddenBitIsOne()._Started.0\ <= false;
                            \Unum::ExponentValueWithBias().0.return.0\ := \Unum::ExponentValueWithBias().0.Unum::HiddenBitIsOne().return.0\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::ExponentValueWithBias().0._State_5\ and ends in state \Unum::ExponentValueWithBias().0._State_5\.
                            --     * The false branch starts in state \Unum::ExponentValueWithBias().0._State_6\ and ends in state \Unum::ExponentValueWithBias().0._State_6\.
                            --     * Execution after either branch will continue in the following state: \Unum::ExponentValueWithBias().0._State_4\.

                            if (\Unum::ExponentValueWithBias().0.return.0\) then 
                                \Unum::ExponentValueWithBias().0._State\ := \Unum::ExponentValueWithBias().0._State_5\;
                            else 
                                \Unum::ExponentValueWithBias().0._State\ := \Unum::ExponentValueWithBias().0._State_6\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentValueWithBias().0._State_4\ => 
                        -- State after the if-else which was started in state \Unum::ExponentValueWithBias().0._State_3\.
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::Exponent()
                        \Unum::ExponentValueWithBias().0.Unum::Exponent()._Started.0\ <= true;
                        \Unum::ExponentValueWithBias().0._State\ := \Unum::ExponentValueWithBias().0._State_7\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentValueWithBias().0._State_5\ => 
                        -- True branch of the if-else started in state \Unum::ExponentValueWithBias().0._State_3\.
                        \Unum::ExponentValueWithBias().0.conditional45e7bd3495aef0adb29743d60986bee4963f49e22dbfea77daec45939a162bd1\ := to_unsigned(0, 32);
                        -- Going to the state after the if-else which was started in state \Unum::ExponentValueWithBias().0._State_3\.
                        if (\Unum::ExponentValueWithBias().0._State\ = \Unum::ExponentValueWithBias().0._State_5\) then 
                            \Unum::ExponentValueWithBias().0._State\ := \Unum::ExponentValueWithBias().0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentValueWithBias().0._State_6\ => 
                        -- False branch of the if-else started in state \Unum::ExponentValueWithBias().0._State_3\.
                        \Unum::ExponentValueWithBias().0.conditional45e7bd3495aef0adb29743d60986bee4963f49e22dbfea77daec45939a162bd1\ := to_unsigned(1, 32);
                        -- Going to the state after the if-else which was started in state \Unum::ExponentValueWithBias().0._State_3\.
                        if (\Unum::ExponentValueWithBias().0._State\ = \Unum::ExponentValueWithBias().0._State_6\) then 
                            \Unum::ExponentValueWithBias().0._State\ := \Unum::ExponentValueWithBias().0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentValueWithBias().0._State_7\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::Exponent()
                        if (\Unum::ExponentValueWithBias().0.Unum::Exponent()._Started.0\ = \Unum::ExponentValueWithBias().0.Unum::Exponent()._Finished.0\) then 
                            \Unum::ExponentValueWithBias().0.Unum::Exponent()._Started.0\ <= false;
                            \Unum::ExponentValueWithBias().0.return.1\ := \Unum::ExponentValueWithBias().0.Unum::Exponent().return.0\;
                            -- Starting state machine invocation for the following method: System.UInt32 Lombiq.Unum.BitMask::GetLowest32Bits()
                            \Unum::ExponentValueWithBias().0.BitMask::GetLowest32Bits().this.parameter.Out.0\ <= \Unum::ExponentValueWithBias().0.return.1\;
                            \Unum::ExponentValueWithBias().0.BitMask::GetLowest32Bits()._Started.0\ <= true;
                            \Unum::ExponentValueWithBias().0._State\ := \Unum::ExponentValueWithBias().0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentValueWithBias().0._State_8\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt32 Lombiq.Unum.BitMask::GetLowest32Bits()
                        if (\Unum::ExponentValueWithBias().0.BitMask::GetLowest32Bits()._Started.0\ = \Unum::ExponentValueWithBias().0.BitMask::GetLowest32Bits()._Finished.0\) then 
                            \Unum::ExponentValueWithBias().0.BitMask::GetLowest32Bits()._Started.0\ <= false;
                            \Unum::ExponentValueWithBias().0.return.2\ := \Unum::ExponentValueWithBias().0.BitMask::GetLowest32Bits().return.0\;
                            -- Starting state machine invocation for the following method: System.Int32 Lombiq.Unum.Unum::Bias()
                            \Unum::ExponentValueWithBias().0.Unum::Bias()._Started.0\ <= true;
                            \Unum::ExponentValueWithBias().0._State\ := \Unum::ExponentValueWithBias().0._State_9\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentValueWithBias().0._State_9\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Int32 Lombiq.Unum.Unum::Bias()
                        if (\Unum::ExponentValueWithBias().0.Unum::Bias()._Started.0\ = \Unum::ExponentValueWithBias().0.Unum::Bias()._Finished.0\) then 
                            \Unum::ExponentValueWithBias().0.Unum::Bias()._Started.0\ <= false;
                            \Unum::ExponentValueWithBias().0.return.3\ := \Unum::ExponentValueWithBias().0.Unum::Bias().return.0\;
                            \Unum::ExponentValueWithBias().0.binaryOperationResult.0\ := \Unum::ExponentValueWithBias().0.return.2\ - unsigned(\Unum::ExponentValueWithBias().0.return.3\);
                            \Unum::ExponentValueWithBias().0.binaryOperationResult.1\ := resize(signed(\Unum::ExponentValueWithBias().0.binaryOperationResult.0\ + \Unum::ExponentValueWithBias().0.conditional45e7bd3495aef0adb29743d60986bee4963f49e22dbfea77daec45939a162bd1\), 32);
                            \Unum::ExponentValueWithBias().0.return\ <= (\Unum::ExponentValueWithBias().0.binaryOperationResult.1\);
                            \Unum::ExponentValueWithBias().0._State\ := \Unum::ExponentValueWithBias().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                end case;
            end if;
        end if;
    end process;
    -- System.Int32 Lombiq.Unum.Unum::ExponentValueWithBias().0 state machine end


    -- System.Boolean Lombiq.Unum.Unum::IsNan().0 state machine start
    \Unum::IsNan().0._StateMachine\: process (\Clock\) 
        Variable \Unum::IsNan().0._State\: \Unum::IsNan().0._States\ := \Unum::IsNan().0._State_0\;
        Variable \Unum::IsNan().0.this\: \Lombiq.Unum.Unum\;
        Variable \Unum::IsNan().0.return.0\: \Lombiq.Unum.BitMask\;
        Variable \Unum::IsNan().0.return.1\: boolean := false;
        Variable \Unum::IsNan().0.return.2\: \Lombiq.Unum.BitMask\;
        Variable \Unum::IsNan().0.return.3\: boolean := false;
        Variable \Unum::IsNan().0.binaryOperationResult.0\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::IsNan().0._Finished\ <= false;
                \Unum::IsNan().0.return\ <= false;
                \Unum::IsNan().0.Unum::get_SignalingNotANumber()._Started.0\ <= false;
                \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ <= false;
                \Unum::IsNan().0.Unum::get_QuietNotANumber()._Started.0\ <= false;
                \Unum::IsNan().0._State\ := \Unum::IsNan().0._State_0\;
                \Unum::IsNan().0.return.1\ := false;
                \Unum::IsNan().0.return.3\ := false;
                \Unum::IsNan().0.binaryOperationResult.0\ := false;
            else 
                case \Unum::IsNan().0._State\ is 
                    when \Unum::IsNan().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::IsNan().0._Started\ = true) then 
                            \Unum::IsNan().0._State\ := \Unum::IsNan().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsNan().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::IsNan().0._Started\ = true) then 
                            \Unum::IsNan().0._Finished\ <= true;
                        else 
                            \Unum::IsNan().0._Finished\ <= false;
                            \Unum::IsNan().0._State\ := \Unum::IsNan().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsNan().0._State_2\ => 
                        \Unum::IsNan().0.this\ := \Unum::IsNan().0.this.parameter.In\;
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_SignalingNotANumber()
                        \Unum::IsNan().0.Unum::get_SignalingNotANumber().this.parameter.Out.0\ <= \Unum::IsNan().0.this\;
                        \Unum::IsNan().0.Unum::get_SignalingNotANumber()._Started.0\ <= true;
                        \Unum::IsNan().0._State\ := \Unum::IsNan().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsNan().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_SignalingNotANumber()
                        if (\Unum::IsNan().0.Unum::get_SignalingNotANumber()._Started.0\ = \Unum::IsNan().0.Unum::get_SignalingNotANumber()._Finished.0\) then 
                            \Unum::IsNan().0.Unum::get_SignalingNotANumber()._Started.0\ <= false;
                            \Unum::IsNan().0.return.0\ := \Unum::IsNan().0.Unum::get_SignalingNotANumber().return.0\;
                            -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.BitMask::op_Equality(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask).left.parameter.Out.0\ <= \Unum::IsNan().0.this\.\UnumBits\;
                            \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask).right.parameter.Out.0\ <= \Unum::IsNan().0.return.0\;
                            \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ <= true;
                            \Unum::IsNan().0._State\ := \Unum::IsNan().0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsNan().0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.BitMask::op_Equality(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ = \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\) then 
                            \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ <= false;
                            \Unum::IsNan().0.return.1\ := \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask).return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_QuietNotANumber()
                            \Unum::IsNan().0.Unum::get_QuietNotANumber().this.parameter.Out.0\ <= \Unum::IsNan().0.this\;
                            \Unum::IsNan().0.Unum::get_QuietNotANumber()._Started.0\ <= true;
                            \Unum::IsNan().0._State\ := \Unum::IsNan().0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsNan().0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_QuietNotANumber()
                        if (\Unum::IsNan().0.Unum::get_QuietNotANumber()._Started.0\ = \Unum::IsNan().0.Unum::get_QuietNotANumber()._Finished.0\) then 
                            \Unum::IsNan().0.Unum::get_QuietNotANumber()._Started.0\ <= false;
                            \Unum::IsNan().0.return.2\ := \Unum::IsNan().0.Unum::get_QuietNotANumber().return.0\;
                            -- The last invocation for the target state machine finished in the previous state, so need to start the next one in the next state.
                            \Unum::IsNan().0._State\ := \Unum::IsNan().0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsNan().0._State_6\ => 
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.BitMask::op_Equality(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask).left.parameter.Out.0\ <= \Unum::IsNan().0.this\.\UnumBits\;
                        \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask).right.parameter.Out.0\ <= \Unum::IsNan().0.return.2\;
                        \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ <= true;
                        \Unum::IsNan().0._State\ := \Unum::IsNan().0._State_7\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsNan().0._State_7\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.BitMask::op_Equality(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ = \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\) then 
                            \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ <= false;
                            \Unum::IsNan().0.return.3\ := \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask).return.0\;
                            \Unum::IsNan().0.binaryOperationResult.0\ := \Unum::IsNan().0.return.1\ or \Unum::IsNan().0.return.3\;
                            \Unum::IsNan().0.return\ <= \Unum::IsNan().0.binaryOperationResult.0\;
                            \Unum::IsNan().0._State\ := \Unum::IsNan().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Lombiq.Unum.Unum::IsNan().0 state machine end


    -- System.Boolean Lombiq.Unum.Unum::IsPositiveInfinity().0 state machine start
    \Unum::IsPositiveInfinity().0._StateMachine\: process (\Clock\) 
        Variable \Unum::IsPositiveInfinity().0._State\: \Unum::IsPositiveInfinity().0._States\ := \Unum::IsPositiveInfinity().0._State_0\;
        Variable \Unum::IsPositiveInfinity().0.this\: \Lombiq.Unum.Unum\;
        Variable \Unum::IsPositiveInfinity().0.return.0\: \Lombiq.Unum.BitMask\;
        Variable \Unum::IsPositiveInfinity().0.return.1\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::IsPositiveInfinity().0._Finished\ <= false;
                \Unum::IsPositiveInfinity().0.return\ <= false;
                \Unum::IsPositiveInfinity().0.Unum::get_PositiveInfinity()._Started.0\ <= false;
                \Unum::IsPositiveInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ <= false;
                \Unum::IsPositiveInfinity().0._State\ := \Unum::IsPositiveInfinity().0._State_0\;
                \Unum::IsPositiveInfinity().0.return.1\ := false;
            else 
                case \Unum::IsPositiveInfinity().0._State\ is 
                    when \Unum::IsPositiveInfinity().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::IsPositiveInfinity().0._Started\ = true) then 
                            \Unum::IsPositiveInfinity().0._State\ := \Unum::IsPositiveInfinity().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsPositiveInfinity().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::IsPositiveInfinity().0._Started\ = true) then 
                            \Unum::IsPositiveInfinity().0._Finished\ <= true;
                        else 
                            \Unum::IsPositiveInfinity().0._Finished\ <= false;
                            \Unum::IsPositiveInfinity().0._State\ := \Unum::IsPositiveInfinity().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsPositiveInfinity().0._State_2\ => 
                        \Unum::IsPositiveInfinity().0.this\ := \Unum::IsPositiveInfinity().0.this.parameter.In\;
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_PositiveInfinity()
                        \Unum::IsPositiveInfinity().0.Unum::get_PositiveInfinity().this.parameter.Out.0\ <= \Unum::IsPositiveInfinity().0.this\;
                        \Unum::IsPositiveInfinity().0.Unum::get_PositiveInfinity()._Started.0\ <= true;
                        \Unum::IsPositiveInfinity().0._State\ := \Unum::IsPositiveInfinity().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsPositiveInfinity().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_PositiveInfinity()
                        if (\Unum::IsPositiveInfinity().0.Unum::get_PositiveInfinity()._Started.0\ = \Unum::IsPositiveInfinity().0.Unum::get_PositiveInfinity()._Finished.0\) then 
                            \Unum::IsPositiveInfinity().0.Unum::get_PositiveInfinity()._Started.0\ <= false;
                            \Unum::IsPositiveInfinity().0.return.0\ := \Unum::IsPositiveInfinity().0.Unum::get_PositiveInfinity().return.0\;
                            -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.BitMask::op_Equality(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \Unum::IsPositiveInfinity().0.BitMask::op_Equality(BitMask,BitMask).left.parameter.Out.0\ <= \Unum::IsPositiveInfinity().0.this\.\UnumBits\;
                            \Unum::IsPositiveInfinity().0.BitMask::op_Equality(BitMask,BitMask).right.parameter.Out.0\ <= \Unum::IsPositiveInfinity().0.return.0\;
                            \Unum::IsPositiveInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ <= true;
                            \Unum::IsPositiveInfinity().0._State\ := \Unum::IsPositiveInfinity().0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsPositiveInfinity().0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.BitMask::op_Equality(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\Unum::IsPositiveInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ = \Unum::IsPositiveInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\) then 
                            \Unum::IsPositiveInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ <= false;
                            \Unum::IsPositiveInfinity().0.return.1\ := \Unum::IsPositiveInfinity().0.BitMask::op_Equality(BitMask,BitMask).return.0\;
                            \Unum::IsPositiveInfinity().0.return\ <= \Unum::IsPositiveInfinity().0.return.1\;
                            \Unum::IsPositiveInfinity().0._State\ := \Unum::IsPositiveInfinity().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Lombiq.Unum.Unum::IsPositiveInfinity().0 state machine end


    -- System.Boolean Lombiq.Unum.Unum::IsNegativeInfinity().0 state machine start
    \Unum::IsNegativeInfinity().0._StateMachine\: process (\Clock\) 
        Variable \Unum::IsNegativeInfinity().0._State\: \Unum::IsNegativeInfinity().0._States\ := \Unum::IsNegativeInfinity().0._State_0\;
        Variable \Unum::IsNegativeInfinity().0.this\: \Lombiq.Unum.Unum\;
        Variable \Unum::IsNegativeInfinity().0.return.0\: \Lombiq.Unum.BitMask\;
        Variable \Unum::IsNegativeInfinity().0.return.1\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::IsNegativeInfinity().0._Finished\ <= false;
                \Unum::IsNegativeInfinity().0.return\ <= false;
                \Unum::IsNegativeInfinity().0.Unum::get_NegativeInfinity()._Started.0\ <= false;
                \Unum::IsNegativeInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ <= false;
                \Unum::IsNegativeInfinity().0._State\ := \Unum::IsNegativeInfinity().0._State_0\;
                \Unum::IsNegativeInfinity().0.return.1\ := false;
            else 
                case \Unum::IsNegativeInfinity().0._State\ is 
                    when \Unum::IsNegativeInfinity().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::IsNegativeInfinity().0._Started\ = true) then 
                            \Unum::IsNegativeInfinity().0._State\ := \Unum::IsNegativeInfinity().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsNegativeInfinity().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::IsNegativeInfinity().0._Started\ = true) then 
                            \Unum::IsNegativeInfinity().0._Finished\ <= true;
                        else 
                            \Unum::IsNegativeInfinity().0._Finished\ <= false;
                            \Unum::IsNegativeInfinity().0._State\ := \Unum::IsNegativeInfinity().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsNegativeInfinity().0._State_2\ => 
                        \Unum::IsNegativeInfinity().0.this\ := \Unum::IsNegativeInfinity().0.this.parameter.In\;
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_NegativeInfinity()
                        \Unum::IsNegativeInfinity().0.Unum::get_NegativeInfinity().this.parameter.Out.0\ <= \Unum::IsNegativeInfinity().0.this\;
                        \Unum::IsNegativeInfinity().0.Unum::get_NegativeInfinity()._Started.0\ <= true;
                        \Unum::IsNegativeInfinity().0._State\ := \Unum::IsNegativeInfinity().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsNegativeInfinity().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_NegativeInfinity()
                        if (\Unum::IsNegativeInfinity().0.Unum::get_NegativeInfinity()._Started.0\ = \Unum::IsNegativeInfinity().0.Unum::get_NegativeInfinity()._Finished.0\) then 
                            \Unum::IsNegativeInfinity().0.Unum::get_NegativeInfinity()._Started.0\ <= false;
                            \Unum::IsNegativeInfinity().0.return.0\ := \Unum::IsNegativeInfinity().0.Unum::get_NegativeInfinity().return.0\;
                            -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.BitMask::op_Equality(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \Unum::IsNegativeInfinity().0.BitMask::op_Equality(BitMask,BitMask).left.parameter.Out.0\ <= \Unum::IsNegativeInfinity().0.this\.\UnumBits\;
                            \Unum::IsNegativeInfinity().0.BitMask::op_Equality(BitMask,BitMask).right.parameter.Out.0\ <= \Unum::IsNegativeInfinity().0.return.0\;
                            \Unum::IsNegativeInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ <= true;
                            \Unum::IsNegativeInfinity().0._State\ := \Unum::IsNegativeInfinity().0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::IsNegativeInfinity().0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.BitMask::op_Equality(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\Unum::IsNegativeInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ = \Unum::IsNegativeInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\) then 
                            \Unum::IsNegativeInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ <= false;
                            \Unum::IsNegativeInfinity().0.return.1\ := \Unum::IsNegativeInfinity().0.BitMask::op_Equality(BitMask,BitMask).return.0\;
                            \Unum::IsNegativeInfinity().0.return\ <= \Unum::IsNegativeInfinity().0.return.1\;
                            \Unum::IsNegativeInfinity().0._State\ := \Unum::IsNegativeInfinity().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Lombiq.Unum.Unum::IsNegativeInfinity().0 state machine end


    -- Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0 state machine start
    \Unum::AddExactUnums(Unum,Unum).0._StateMachine\: process (\Clock\) 
        Variable \Unum::AddExactUnums(Unum,Unum).0._State\: \Unum::AddExactUnums(Unum,Unum).0._States\ := \Unum::AddExactUnums(Unum,Unum).0._State_0\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.left\: \Lombiq.Unum.Unum\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.right\: \Lombiq.Unum.Unum\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.bitMask\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.flag\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.result\: \Lombiq.Unum.Unum\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.flag2\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.flag3\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.flag4\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.unum\: \Lombiq.Unum.Unum\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.num\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::AddExactUnums(Unum,Unum).0.flag5\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.flag6\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.num2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::AddExactUnums(Unum,Unum).0.right2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::AddExactUnums(Unum,Unum).0.num3\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::AddExactUnums(Unum,Unum).0.flag7\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.flag8\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.signBit\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.flag9\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.num4\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::AddExactUnums(Unum,Unum).0.exponent\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.exponentSize\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Unum::AddExactUnums(Unum,Unum).0.uncertainityBit\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.flag10\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.num5\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.flag11\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.flag12\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.flag13\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.0\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.1\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.0\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.2\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.3\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.4\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.1\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.5\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.6\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.2\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.3\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.7\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.8\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.9\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.4\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.10\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.11\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.12\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.5\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.13\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.14\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.15\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.6\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.16\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.17\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.7\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.8\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.18\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.19\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.9\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.20\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.10\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.11\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.21\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.12\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.22\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.13\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.14\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.23\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.24\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.25\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.26\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.27\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.28\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.29\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.15\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.30\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.31\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.32\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.33\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.34\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.35\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.36\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.37\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.38\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.16\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.39\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.40\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.41\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.17\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.42\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.18\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.19\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.43\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.20\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.44\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.21\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.22\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.23\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.45\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.46\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.47\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.48\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.49\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.50\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.51\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.52\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.24\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.53\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.25\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.26\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.54\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.27\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.55\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.28\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.29\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.30\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.56\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.57\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.58\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.59\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.60\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.61\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.62\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.31\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.32\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::AddExactUnums(Unum,Unum).0.objectb27a734c21885631ebb68e1234fb9c8390b7e1444b1d60f27d01ade0c7b5d9bc\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.33\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.63\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.64\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.65\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.34\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.66\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.67\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.35\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.68\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.36\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.69\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.37\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.70\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.38\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.71\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.39\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.40\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.72\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.73\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.41\: boolean := false;
        Variable \Unum::AddExactUnums(Unum,Unum).0.return.74\: \Lombiq.Unum.BitMask\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::AddExactUnums(Unum,Unum).0._Finished\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNan()._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber()._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask)._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity()._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity()._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::get_PositiveInfinity()._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::get_NegativeInfinity()._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment)._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\ <= to_signed(0, 32);
                \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean).signBitsMatch.parameter.Out.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean)._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne()._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction()._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_GreaterThanOrEqual(BitMask,BitMask)._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::get_Size()._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueToExponentBits(Int32,Byte).value.parameter.Out.0\ <= to_signed(0, 32);
                \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueToExponentBits(Int32,Byte).size.parameter.Out.0\ <= to_unsigned(0, 8);
                \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueToExponentBits(Int32,Byte)._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.BitMask::ShiftOutLeastSignificantZeros()._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.BitMask::SetZero(UInt16).index.parameter.Out.0\ <= to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.BitMask::SetZero(UInt16)._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::IsExact()._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).signBit.parameter.Out.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).uncertainityBit.parameter.Out.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).exponentSize.parameter.Out.0\ <= to_unsigned(0, 8);
                \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).fractionSize.parameter.Out.0\ <= to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Started.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_0\;
                \Unum::AddExactUnums(Unum,Unum).0.flag\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.flag2\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.flag3\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.flag4\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.num\ := to_signed(0, 32);
                \Unum::AddExactUnums(Unum,Unum).0.flag5\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.flag6\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.num2\ := to_signed(0, 32);
                \Unum::AddExactUnums(Unum,Unum).0.right2\ := to_signed(0, 32);
                \Unum::AddExactUnums(Unum,Unum).0.num3\ := to_signed(0, 32);
                \Unum::AddExactUnums(Unum,Unum).0.flag7\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.flag8\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.signBit\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.flag9\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.num4\ := to_signed(0, 32);
                \Unum::AddExactUnums(Unum,Unum).0.exponentSize\ := to_unsigned(0, 8);
                \Unum::AddExactUnums(Unum,Unum).0.uncertainityBit\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.flag10\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.num5\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.flag11\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.flag12\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.flag13\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.0\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.1\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.0\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.3\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.4\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.1\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.5\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.6\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.2\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.3\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.8\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.9\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.4\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.11\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.12\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.5\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.14\ := to_signed(0, 32);
                \Unum::AddExactUnums(Unum,Unum).0.return.15\ := to_signed(0, 32);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.6\ := to_signed(0, 32);
                \Unum::AddExactUnums(Unum,Unum).0.return.16\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.17\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.7\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.8\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.18\ := to_signed(0, 32);
                \Unum::AddExactUnums(Unum,Unum).0.return.19\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.9\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.return.20\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.10\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.11\ := to_signed(0, 32);
                \Unum::AddExactUnums(Unum,Unum).0.return.21\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.12\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.return.22\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.13\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.14\ := to_signed(0, 32);
                \Unum::AddExactUnums(Unum,Unum).0.return.28\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.29\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.15\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.32\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.33\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.34\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.35\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.36\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.37\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.38\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.16\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.39\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.40\ := to_signed(0, 32);
                \Unum::AddExactUnums(Unum,Unum).0.return.41\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.17\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.return.42\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.18\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.19\ := to_signed(0, 32);
                \Unum::AddExactUnums(Unum,Unum).0.return.43\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.20\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.return.44\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.21\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.22\ := to_signed(0, 32);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.23\ := to_signed(0, 32);
                \Unum::AddExactUnums(Unum,Unum).0.return.50\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.51\ := to_signed(0, 32);
                \Unum::AddExactUnums(Unum,Unum).0.return.52\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.24\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.return.53\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.25\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.26\ := to_signed(0, 32);
                \Unum::AddExactUnums(Unum,Unum).0.return.54\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.27\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.return.55\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.28\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.29\ := to_signed(0, 32);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.30\ := to_signed(0, 32);
                \Unum::AddExactUnums(Unum,Unum).0.return.61\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.return.62\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.31\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.32\ := to_signed(0, 32);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.33\ := to_signed(0, 32);
                \Unum::AddExactUnums(Unum,Unum).0.return.63\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.34\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.67\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.35\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.68\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.36\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.return.69\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.37\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.70\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.38\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.39\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.40\ := to_unsigned(0, 16);
                \Unum::AddExactUnums(Unum,Unum).0.return.72\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.return.73\ := false;
                \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.41\ := false;
            else 
                case \Unum::AddExactUnums(Unum,Unum).0._State\ is 
                    when \Unum::AddExactUnums(Unum,Unum).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::AddExactUnums(Unum,Unum).0._Started\ = true) then 
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::AddExactUnums(Unum,Unum).0._Started\ = true) then 
                            \Unum::AddExactUnums(Unum,Unum).0._Finished\ <= true;
                        else 
                            \Unum::AddExactUnums(Unum,Unum).0._Finished\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_2\ => 
                        \Unum::AddExactUnums(Unum,Unum).0.left\ := \Unum::AddExactUnums(Unum,Unum).0.left.parameter.In\;
                        \Unum::AddExactUnums(Unum,Unum).0.right\ := \Unum::AddExactUnums(Unum,Unum).0.right.parameter.In\;
                        -- Initializing record fields to their defaults.
                        \Unum::AddExactUnums(Unum,Unum).0.bitMask\.\IsNull\ := false;
                        \Unum::AddExactUnums(Unum,Unum).0.bitMask\.\Size\ := to_unsigned(0, 16);
                        \Unum::AddExactUnums(Unum,Unum).0.bitMask\.\SegmentCount\ := to_unsigned(0, 16);
                        \Unum::AddExactUnums(Unum,Unum).0.bitMask\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                        \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.bitMask\;
                        \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\.\_environment\.\Size\;
                        \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\ <= False;
                        \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.bitMask\ := \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\;
                            -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::IsNan()
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNan().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNan()._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::IsNan()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::IsNan()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNan()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNan()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.0\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNan().return.0\;
                            -- The last invocation for the target state machine just finished, so need to start the next one in a later state.
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_5\ => 
                        -- This state was just added to leave time for the invocation proxy to register that the previous invocation finished.
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_6\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_6\ => 
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::IsNan()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNan().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.right\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNan()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_7\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_7\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::IsNan()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::IsNan()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNan()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNan()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.1\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNan().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.0\ := \Unum::AddExactUnums(Unum,Unum).0.return.0\ or \Unum::AddExactUnums(Unum,Unum).0.return.1\;
                            \Unum::AddExactUnums(Unum,Unum).0.flag\ := \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.0\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_9\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_11\.
                            --     * The false branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_12\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_19\.
                            --     * Execution after either branch will continue in the following state: \Unum::AddExactUnums(Unum,Unum).0._State_8\.

                            if (\Unum::AddExactUnums(Unum,Unum).0.flag\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_9\;
                            else 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_12\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_8\ => 
                        -- State after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_7\.
                        \Unum::AddExactUnums(Unum,Unum).0.return\ <= \Unum::AddExactUnums(Unum,Unum).0.result\;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_9\ => 
                        -- True branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_7\.
                        -- Initializing record fields to their defaults.
                        \Unum::AddExactUnums(Unum,Unum).0.result\.\IsNull\ := false;
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_QuietNotANumber()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_10\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_10\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_QuietNotANumber()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.2\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber().return.0\;
                            -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,Lombiq.Unum.BitMask)
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.result\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).environment.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\.\_environment\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).bits.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.return.2\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask)._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_11\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_11\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,Lombiq.Unum.BitMask)
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask)._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask)._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask)._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.result\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).this.parameter.In.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.left\.\_environment\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).environment.parameter.In.0\;
                            -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_7\.
                            if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_11\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_8\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_12\ => 
                        -- False branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_7\.
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::IsPositiveInfinity()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_13\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_13\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::IsPositiveInfinity()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.3\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity().return.0\;
                            -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::IsNegativeInfinity()
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.right\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity()._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_14\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_14\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::IsNegativeInfinity()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.4\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.1\ := \Unum::AddExactUnums(Unum,Unum).0.return.3\ and \Unum::AddExactUnums(Unum,Unum).0.return.4\;
                            -- The last invocation for the target state machine just finished, so need to start the next one in a later state.
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_15\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_15\ => 
                        -- This state was just added to leave time for the invocation proxy to register that the previous invocation finished.
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_16\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_16\ => 
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::IsNegativeInfinity()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_17\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_17\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::IsNegativeInfinity()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.5\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity().return.0\;
                            -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::IsPositiveInfinity()
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.right\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity()._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_18\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_18\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::IsPositiveInfinity()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.6\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.2\ := \Unum::AddExactUnums(Unum,Unum).0.return.5\ and \Unum::AddExactUnums(Unum,Unum).0.return.6\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.3\ := \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.1\ or \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.2\;
                            \Unum::AddExactUnums(Unum,Unum).0.flag2\ := \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.3\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_20\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_22\.
                            --     * The false branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_23\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_28\.
                            --     * Execution after either branch will continue in the following state: \Unum::AddExactUnums(Unum,Unum).0._State_19\.

                            if (\Unum::AddExactUnums(Unum,Unum).0.flag2\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_20\;
                            else 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_23\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \Unum::AddExactUnums(Unum,Unum).0._State_19\ => 
                        -- State after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_18\.
                        -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_7\.
                        if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_19\) then 
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_20\ => 
                        -- True branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_18\.
                        -- Initializing record fields to their defaults.
                        \Unum::AddExactUnums(Unum,Unum).0.result\.\IsNull\ := false;
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_QuietNotANumber()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_21\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_21\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_QuietNotANumber()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.7\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber().return.0\;
                            -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,Lombiq.Unum.BitMask)
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.result\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).environment.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\.\_environment\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).bits.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.return.7\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask)._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_22\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_22\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,Lombiq.Unum.BitMask)
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask)._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask)._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask)._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.result\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).this.parameter.In.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.left\.\_environment\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).environment.parameter.In.0\;
                            -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_18\.
                            if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_22\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_19\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_23\ => 
                        -- False branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_18\.
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::IsPositiveInfinity()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_24\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_24\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::IsPositiveInfinity()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.8\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity().return.0\;
                            -- The last invocation for the target state machine just finished, so need to start the next one in a later state.
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_25\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_25\ => 
                        -- This state was just added to leave time for the invocation proxy to register that the previous invocation finished.
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_26\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_26\ => 
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::IsPositiveInfinity()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.right\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_27\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_27\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::IsPositiveInfinity()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.9\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.4\ := \Unum::AddExactUnums(Unum,Unum).0.return.8\ or \Unum::AddExactUnums(Unum,Unum).0.return.9\;
                            \Unum::AddExactUnums(Unum,Unum).0.flag3\ := \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.4\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_29\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_31\.
                            --     * The false branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_32\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_37\.
                            --     * Execution after either branch will continue in the following state: \Unum::AddExactUnums(Unum,Unum).0._State_28\.

                            if (\Unum::AddExactUnums(Unum,Unum).0.flag3\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_29\;
                            else 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_32\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_28\ => 
                        -- State after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_27\.
                        -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_18\.
                        if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_28\) then 
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_19\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_29\ => 
                        -- True branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_27\.
                        -- Initializing record fields to their defaults.
                        \Unum::AddExactUnums(Unum,Unum).0.result\.\IsNull\ := false;
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_PositiveInfinity()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::get_PositiveInfinity().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::get_PositiveInfinity()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_30\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_30\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_PositiveInfinity()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::get_PositiveInfinity()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::get_PositiveInfinity()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_PositiveInfinity()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.10\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::get_PositiveInfinity().return.0\;
                            -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,Lombiq.Unum.BitMask)
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.result\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).environment.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\.\_environment\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).bits.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.return.10\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask)._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_31\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_31\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,Lombiq.Unum.BitMask)
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask)._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask)._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask)._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.result\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).this.parameter.In.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.left\.\_environment\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).environment.parameter.In.0\;
                            -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_27\.
                            if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_31\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_28\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_32\ => 
                        -- False branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_27\.
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::IsNegativeInfinity()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_33\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_33\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::IsNegativeInfinity()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.11\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity().return.0\;
                            -- The last invocation for the target state machine just finished, so need to start the next one in a later state.
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_34\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_34\ => 
                        -- This state was just added to leave time for the invocation proxy to register that the previous invocation finished.
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_35\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_35\ => 
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::IsNegativeInfinity()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.right\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_36\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_36\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::IsNegativeInfinity()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.12\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.5\ := \Unum::AddExactUnums(Unum,Unum).0.return.11\ or \Unum::AddExactUnums(Unum,Unum).0.return.12\;
                            \Unum::AddExactUnums(Unum,Unum).0.flag4\ := \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.5\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_38\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_40\.
                            --     * The false branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_41\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_155\.
                            --     * Execution after either branch will continue in the following state: \Unum::AddExactUnums(Unum,Unum).0._State_37\.

                            if (\Unum::AddExactUnums(Unum,Unum).0.flag4\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_38\;
                            else 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_41\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_37\ => 
                        -- State after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_36\.
                        -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_27\.
                        if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_37\) then 
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_28\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_38\ => 
                        -- True branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_36\.
                        -- Initializing record fields to their defaults.
                        \Unum::AddExactUnums(Unum,Unum).0.result\.\IsNull\ := false;
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_NegativeInfinity()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::get_NegativeInfinity().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::get_NegativeInfinity()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_39\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_39\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_NegativeInfinity()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::get_NegativeInfinity()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::get_NegativeInfinity()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_NegativeInfinity()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.13\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::get_NegativeInfinity().return.0\;
                            -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,Lombiq.Unum.BitMask)
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.result\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).environment.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\.\_environment\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).bits.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.return.13\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask)._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_40\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_40\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,Lombiq.Unum.BitMask)
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask)._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask)._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask)._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.result\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).this.parameter.In.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.left\.\_environment\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).environment.parameter.In.0\;
                            -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_36\.
                            if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_40\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_37\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_41\ => 
                        -- False branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_36\.
                        -- Initializing record fields to their defaults.
                        \Unum::AddExactUnums(Unum,Unum).0.unum\.\IsNull\ := false;
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment)
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment).this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.unum\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment).environment.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\.\_environment\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment)._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_42\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_42\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment)
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment)._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment)._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment)._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.unum\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment).this.parameter.In.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.left\.\_environment\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment).environment.parameter.In.0\;
                            -- Starting state machine invocation for the following method: System.Int32 Lombiq.Unum.Unum::ExponentValueWithBias()
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_43\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_43\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Int32 Lombiq.Unum.Unum::ExponentValueWithBias()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.14\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias().return.0\;
                            -- The last invocation for the target state machine just finished, so need to start the next one in a later state.
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_44\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_44\ => 
                        -- This state was just added to leave time for the invocation proxy to register that the previous invocation finished.
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_45\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_45\ => 
                        -- Starting state machine invocation for the following method: System.Int32 Lombiq.Unum.Unum::ExponentValueWithBias()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.right\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_46\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_46\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Int32 Lombiq.Unum.Unum::ExponentValueWithBias()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.15\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.6\ := \Unum::AddExactUnums(Unum,Unum).0.return.14\ - \Unum::AddExactUnums(Unum,Unum).0.return.15\;
                            \Unum::AddExactUnums(Unum,Unum).0.num\ := \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.6\;
                            -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::IsPositive()
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_47\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_47\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::IsPositive()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.16\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive().return.0\;
                            -- The last invocation for the target state machine just finished, so need to start the next one in a later state.
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_48\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_48\ => 
                        -- This state was just added to leave time for the invocation proxy to register that the previous invocation finished.
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_49\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_49\ => 
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::IsPositive()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.right\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_50\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_50\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::IsPositive()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.17\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.7\ := \Unum::AddExactUnums(Unum,Unum).0.return.16\ = \Unum::AddExactUnums(Unum,Unum).0.return.17\;
                            \Unum::AddExactUnums(Unum,Unum).0.flag5\ := \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.7\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.8\ := \Unum::AddExactUnums(Unum,Unum).0.num\ = to_signed(0, 32);
                            \Unum::AddExactUnums(Unum,Unum).0.flag6\ := \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.8\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_52\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_65\.
                            --     * The false branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_95\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_96\.
                            --     * Execution after either branch will continue in the following state: \Unum::AddExactUnums(Unum,Unum).0._State_51\.

                            if (\Unum::AddExactUnums(Unum,Unum).0.flag6\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_52\;
                            else 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_95\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \Unum::AddExactUnums(Unum,Unum).0._State_51\ => 
                        -- State after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_50\.
                        -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.BitMask::GetMostSignificantOnePosition()
                        \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.bitMask\;
                        \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_125\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_52\ => 
                        -- True branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_50\.
                        -- Starting state machine invocation for the following method: System.Int32 Lombiq.Unum.Unum::ExponentValueWithBias()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_53\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_53\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Int32 Lombiq.Unum.Unum::ExponentValueWithBias()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.18\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.num2\ := \Unum::AddExactUnums(Unum,Unum).0.return.18\;
                            -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::get_FractionSizeMax()
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.unum\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_54\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_54\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::get_FractionSizeMax()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.19\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.9\ := \Unum::AddExactUnums(Unum,Unum).0.return.19\ + to_unsigned(1, 16);
                            -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::FractionSize()
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_55\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_55\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::FractionSize()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.20\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.10\ := \Unum::AddExactUnums(Unum,Unum).0.return.20\ + to_unsigned(1, 16);
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.11\ := resize(signed(\Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.9\ - \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.10\), 32);
                            \Unum::AddExactUnums(Unum,Unum).0.right2\ := (\Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.11\);
                            -- The last invocation for the target state machine finished in the previous state, so need to start the next one in the next state.
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_56\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \Unum::AddExactUnums(Unum,Unum).0._State_56\ => 
                        -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::get_FractionSizeMax()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.unum\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_57\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_57\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::get_FractionSizeMax()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.21\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.12\ := \Unum::AddExactUnums(Unum,Unum).0.return.21\ + to_unsigned(1, 16);
                            -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::FractionSize()
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.right\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_58\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_58\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::FractionSize()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.22\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.13\ := \Unum::AddExactUnums(Unum,Unum).0.return.22\ + to_unsigned(1, 16);
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.14\ := resize(signed(\Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.12\ - \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.13\), 32);
                            \Unum::AddExactUnums(Unum,Unum).0.num3\ := (\Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.14\);
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit()
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_59\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \Unum::AddExactUnums(Unum,Unum).0._State_59\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.23\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit().return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.return.23\;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.right2\;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_60\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_60\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.24\ := \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).return.0\;
                            -- The last invocation for the target state machine finished in the previous state, so need to start the next one in the next state.
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_61\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_61\ => 
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.right\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_62\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_62\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.25\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit().return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.return.25\;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.num3\;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_63\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_63\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.26\ := \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::AddAlignedFractions(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean)
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean).left.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.return.24\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean).right.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.return.26\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean).signBitsMatch.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.flag5\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean)._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_64\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_64\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::AddAlignedFractions(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean)
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean)._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean)._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean)._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.27\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean).return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.bitMask\ := \Unum::AddExactUnums(Unum,Unum).0.return.27\;
                            \Unum::AddExactUnums(Unum,Unum).0.flag7\ := not(\Unum::AddExactUnums(Unum,Unum).0.flag5\);

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_66\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_71\.
                            --     * The false branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_92\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_94\.
                            --     * Execution after either branch will continue in the following state: \Unum::AddExactUnums(Unum,Unum).0._State_65\.

                            if (\Unum::AddExactUnums(Unum,Unum).0.flag7\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_66\;
                            else 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_92\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_65\ => 
                        -- State after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_64\.
                        -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_50\.
                        if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_65\) then 
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_51\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_66\ => 
                        -- True branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_64\.
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::HiddenBitIsOne()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_67\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_67\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::HiddenBitIsOne()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.28\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne().return.0\;
                            -- The last invocation for the target state machine just finished, so need to start the next one in a later state.
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_68\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_68\ => 
                        -- This state was just added to leave time for the invocation proxy to register that the previous invocation finished.
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_69\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_69\ => 
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::HiddenBitIsOne()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.right\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_70\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_70\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::HiddenBitIsOne()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.29\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.15\ := \Unum::AddExactUnums(Unum,Unum).0.return.28\ = \Unum::AddExactUnums(Unum,Unum).0.return.29\;
                            \Unum::AddExactUnums(Unum,Unum).0.flag8\ := \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.15\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_72\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_78\.
                            --     * The false branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_84\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_86\.
                            --     * Execution after either branch will continue in the following state: \Unum::AddExactUnums(Unum,Unum).0._State_71\.

                            if (\Unum::AddExactUnums(Unum,Unum).0.flag8\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_72\;
                            else 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_84\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_71\ => 
                        -- State after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_70\.
                        -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_64\.
                        if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_71\) then 
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_65\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_72\ => 
                        -- True branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_70\.
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::Fraction()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_73\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_73\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::Fraction()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.30\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction().return.0\;
                            -- The last invocation for the target state machine just finished, so need to start the next one in a later state.
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_74\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_74\ => 
                        -- This state was just added to leave time for the invocation proxy to register that the previous invocation finished.
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_75\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_75\ => 
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::Fraction()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.right\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_76\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_76\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::Fraction()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.31\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction().return.0\;
                            -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.BitMask::op_GreaterThanOrEqual(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_GreaterThanOrEqual(BitMask,BitMask).left.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.return.30\;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_GreaterThanOrEqual(BitMask,BitMask).right.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.return.31\;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_GreaterThanOrEqual(BitMask,BitMask)._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_77\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_77\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.BitMask::op_GreaterThanOrEqual(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::op_GreaterThanOrEqual(BitMask,BitMask)._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_GreaterThanOrEqual(BitMask,BitMask)._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_GreaterThanOrEqual(BitMask,BitMask)._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.32\ := \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_GreaterThanOrEqual(BitMask,BitMask).return.0\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_79\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_80\.
                            --     * The false branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_81\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_83\.
                            --     * Execution after either branch will continue in the following state: \Unum::AddExactUnums(Unum,Unum).0._State_78\.

                            if (\Unum::AddExactUnums(Unum,Unum).0.return.32\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_79\;
                            else 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_81\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_78\ => 
                        -- State after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_77\.
                        -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_70\.
                        if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_78\) then 
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_71\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_79\ => 
                        -- True branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_77\.
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::IsPositive()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_80\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_80\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::IsPositive()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.33\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.signBit\ := not(\Unum::AddExactUnums(Unum,Unum).0.return.33\);
                            -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_77\.
                            if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_80\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_78\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_81\ => 
                        -- False branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_77\.
                        -- The last invocation for the target state machine finished in the previous state, so need to start the next one in the next state.
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_82\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_82\ => 
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::IsPositive()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.right\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_83\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_83\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::IsPositive()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.34\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.signBit\ := not(\Unum::AddExactUnums(Unum,Unum).0.return.34\);
                            -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_77\.
                            if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_83\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_78\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_84\ => 
                        -- False branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_70\.
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::HiddenBitIsOne()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_85\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_85\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::HiddenBitIsOne()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.35\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne().return.0\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_87\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_88\.
                            --     * The false branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_89\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_91\.
                            --     * Execution after either branch will continue in the following state: \Unum::AddExactUnums(Unum,Unum).0._State_86\.

                            if (\Unum::AddExactUnums(Unum,Unum).0.return.35\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_87\;
                            else 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_89\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_86\ => 
                        -- State after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_85\.
                        -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_70\.
                        if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_86\) then 
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_71\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_87\ => 
                        -- True branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_85\.
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::IsPositive()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_88\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_88\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::IsPositive()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.36\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.signBit\ := not(\Unum::AddExactUnums(Unum,Unum).0.return.36\);
                            -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_85\.
                            if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_88\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_86\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_89\ => 
                        -- False branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_85\.
                        -- The last invocation for the target state machine finished in the previous state, so need to start the next one in the next state.
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_90\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_90\ => 
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::IsPositive()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.right\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_91\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_91\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::IsPositive()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.37\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.signBit\ := not(\Unum::AddExactUnums(Unum,Unum).0.return.37\);
                            -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_85\.
                            if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_91\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_86\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_92\ => 
                        -- False branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_64\.
                        -- The last invocation for the target state machine finished in the previous state, so need to start the next one in the next state.
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_93\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_93\ => 
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::IsPositive()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_94\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_94\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::IsPositive()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.38\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.signBit\ := not(\Unum::AddExactUnums(Unum,Unum).0.return.38\);
                            -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_64\.
                            if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_94\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_65\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_95\ => 
                        -- False branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_50\.
                        \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.16\ := \Unum::AddExactUnums(Unum,Unum).0.num\ > to_signed(0, 32);
                        \Unum::AddExactUnums(Unum,Unum).0.flag9\ := \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.16\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_97\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_110\.
                        --     * The false branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_111\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_124\.
                        --     * Execution after either branch will continue in the following state: \Unum::AddExactUnums(Unum,Unum).0._State_96\.

                        if (\Unum::AddExactUnums(Unum,Unum).0.flag9\) then 
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_97\;
                        else 
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_111\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_96\ => 
                        -- State after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_95\.
                        -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_50\.
                        if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_96\) then 
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_51\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_97\ => 
                        -- True branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_95\.
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::IsPositive()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_98\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_98\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::IsPositive()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.39\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.signBit\ := not(\Unum::AddExactUnums(Unum,Unum).0.return.39\);
                            -- Starting state machine invocation for the following method: System.Int32 Lombiq.Unum.Unum::ExponentValueWithBias()
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_99\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_99\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Int32 Lombiq.Unum.Unum::ExponentValueWithBias()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.40\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.num2\ := \Unum::AddExactUnums(Unum,Unum).0.return.40\;
                            -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::get_FractionSizeMax()
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.unum\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_100\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_100\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::get_FractionSizeMax()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.41\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.17\ := \Unum::AddExactUnums(Unum,Unum).0.return.41\ + to_unsigned(1, 16);
                            -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::FractionSize()
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_101\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_101\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::FractionSize()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.42\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.18\ := \Unum::AddExactUnums(Unum,Unum).0.return.42\ + to_unsigned(1, 16);
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.19\ := resize(signed(\Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.17\ - \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.18\), 32);
                            \Unum::AddExactUnums(Unum,Unum).0.right2\ := (\Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.19\);
                            -- The last invocation for the target state machine finished in the previous state, so need to start the next one in the next state.
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_102\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \Unum::AddExactUnums(Unum,Unum).0._State_102\ => 
                        -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::get_FractionSizeMax()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.unum\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_103\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_103\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::get_FractionSizeMax()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.43\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.20\ := \Unum::AddExactUnums(Unum,Unum).0.return.43\ + to_unsigned(1, 16);
                            -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::FractionSize()
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.right\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_104\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_104\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::FractionSize()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.44\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.21\ := \Unum::AddExactUnums(Unum,Unum).0.return.44\ + to_unsigned(1, 16);
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.22\ := resize(signed(\Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.20\ - \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.21\), 32);
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.23\ := resize((\Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.22\) - \Unum::AddExactUnums(Unum,Unum).0.num\, 32);
                            \Unum::AddExactUnums(Unum,Unum).0.num3\ := \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.23\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit()
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_105\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \Unum::AddExactUnums(Unum,Unum).0._State_105\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.45\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit().return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.return.45\;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.right2\;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_106\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_106\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.46\ := \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.bitMask\ := \Unum::AddExactUnums(Unum,Unum).0.return.46\;
                            -- The last invocation for the target state machine finished in the previous state, so need to start the next one in the next state.
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_107\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_107\ => 
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.right\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_108\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_108\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.47\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit().return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.return.47\;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.num3\;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_109\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_109\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.48\ := \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::AddAlignedFractions(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean)
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean).left.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.bitMask\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean).right.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.return.48\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean).signBitsMatch.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.flag5\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean)._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_110\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_110\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::AddAlignedFractions(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean)
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean)._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean)._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean)._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.49\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean).return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.bitMask\ := \Unum::AddExactUnums(Unum,Unum).0.return.49\;
                            -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_95\.
                            if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_110\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_96\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_111\ => 
                        -- False branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_95\.
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::IsPositive()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.right\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_112\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_112\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::IsPositive()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.50\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.signBit\ := not(\Unum::AddExactUnums(Unum,Unum).0.return.50\);
                            -- Starting state machine invocation for the following method: System.Int32 Lombiq.Unum.Unum::ExponentValueWithBias()
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.right\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_113\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_113\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Int32 Lombiq.Unum.Unum::ExponentValueWithBias()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.51\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.num2\ := \Unum::AddExactUnums(Unum,Unum).0.return.51\;
                            -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::get_FractionSizeMax()
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.unum\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_114\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_114\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::get_FractionSizeMax()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.52\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.24\ := \Unum::AddExactUnums(Unum,Unum).0.return.52\ + to_unsigned(1, 16);
                            -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::FractionSize()
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.right\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_115\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_115\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::FractionSize()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.53\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.25\ := \Unum::AddExactUnums(Unum,Unum).0.return.53\ + to_unsigned(1, 16);
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.26\ := resize(signed(\Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.24\ - \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.25\), 32);
                            \Unum::AddExactUnums(Unum,Unum).0.right2\ := (\Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.26\);
                            -- The last invocation for the target state machine finished in the previous state, so need to start the next one in the next state.
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_116\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \Unum::AddExactUnums(Unum,Unum).0._State_116\ => 
                        -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::get_FractionSizeMax()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.unum\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_117\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_117\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::get_FractionSizeMax()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.54\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.27\ := \Unum::AddExactUnums(Unum,Unum).0.return.54\ + to_unsigned(1, 16);
                            -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::FractionSize()
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_118\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_118\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::FractionSize()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.55\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.28\ := \Unum::AddExactUnums(Unum,Unum).0.return.55\ + to_unsigned(1, 16);
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.29\ := resize(signed(\Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.27\ - \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.28\), 32);
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.30\ := resize((\Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.29\) + \Unum::AddExactUnums(Unum,Unum).0.num\, 32);
                            \Unum::AddExactUnums(Unum,Unum).0.num3\ := \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.30\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit()
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.right\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_119\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \Unum::AddExactUnums(Unum,Unum).0._State_119\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.56\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit().return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.return.56\;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.right2\;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_120\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_120\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.57\ := \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.bitMask\ := \Unum::AddExactUnums(Unum,Unum).0.return.57\;
                            -- The last invocation for the target state machine finished in the previous state, so need to start the next one in the next state.
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_121\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_121\ => 
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_122\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_122\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.58\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit().return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.return.58\;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.num3\;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_123\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_123\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32)
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.59\ := \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::AddAlignedFractions(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean)
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean).left.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.bitMask\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean).right.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.return.59\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean).signBitsMatch.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.flag5\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean)._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_124\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_124\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::AddAlignedFractions(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean)
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean)._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean)._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean)._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.60\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean).return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.bitMask\ := \Unum::AddExactUnums(Unum,Unum).0.return.60\;
                            -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_95\.
                            if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_124\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_96\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_125\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.BitMask::GetMostSignificantOnePosition()
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.61\ := \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition().return.0\;
                            -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::get_FractionSizeMax()
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.unum\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_126\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_126\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::get_FractionSizeMax()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.62\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.31\ := \Unum::AddExactUnums(Unum,Unum).0.return.62\ + to_unsigned(1, 16);
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.32\ := resize(signed(\Unum::AddExactUnums(Unum,Unum).0.return.61\ - \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.31\), 32);
                            \Unum::AddExactUnums(Unum,Unum).0.num4\ := (\Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.32\);
                            -- Initializing record fields to their defaults.
                            \Unum::AddExactUnums(Unum,Unum).0.objectb27a734c21885631ebb68e1234fb9c8390b7e1444b1d60f27d01ade0c7b5d9bc\.\IsNull\ := false;
                            \Unum::AddExactUnums(Unum,Unum).0.objectb27a734c21885631ebb68e1234fb9c8390b7e1444b1d60f27d01ade0c7b5d9bc\.\Size\ := to_unsigned(0, 16);
                            \Unum::AddExactUnums(Unum,Unum).0.objectb27a734c21885631ebb68e1234fb9c8390b7e1444b1d60f27d01ade0c7b5d9bc\.\SegmentCount\ := to_unsigned(0, 16);
                            \Unum::AddExactUnums(Unum,Unum).0.objectb27a734c21885631ebb68e1234fb9c8390b7e1444b1d60f27d01ade0c7b5d9bc\.\Segments\ := (others => to_unsigned(0, 32));
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.objectb27a734c21885631ebb68e1234fb9c8390b7e1444b1d60f27d01ade0c7b5d9bc\;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\.\_environment\.\Size\;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\ <= False;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_127\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \Unum::AddExactUnums(Unum,Unum).0._State_127\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.objectb27a734c21885631ebb68e1234fb9c8390b7e1444b1d60f27d01ade0c7b5d9bc\ := \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.33\ := \Unum::AddExactUnums(Unum,Unum).0.num2\ + \Unum::AddExactUnums(Unum,Unum).0.num4\;
                            -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.Unum::get_Size()
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_Size().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_Size()._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_128\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_128\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.Unum::get_Size()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::get_Size()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::get_Size()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_Size()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.63\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::get_Size().return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentValueToExponentBits(System.Int32,System.Byte)
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueToExponentBits(Int32,Byte).value.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.33\;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueToExponentBits(Int32,Byte).size.parameter.Out.0\ <= resize(\Unum::AddExactUnums(Unum,Unum).0.return.63\, 8);
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueToExponentBits(Int32,Byte)._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_129\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_129\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentValueToExponentBits(System.Int32,System.Byte)
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueToExponentBits(Int32,Byte)._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueToExponentBits(Int32,Byte)._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueToExponentBits(Int32,Byte)._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.64\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueToExponentBits(Int32,Byte).return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_Addition(BitMask,BitMask).left.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.objectb27a734c21885631ebb68e1234fb9c8390b7e1444b1d60f27d01ade0c7b5d9bc\;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_Addition(BitMask,BitMask).right.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.return.64\;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_130\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_130\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.65\ := \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_Addition(BitMask,BitMask).return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.exponent\ := \Unum::AddExactUnums(Unum,Unum).0.return.65\;
                            \Unum::AddExactUnums(Unum,Unum).0.exponentSize\ := to_unsigned(0, 8);
                            \Unum::AddExactUnums(Unum,Unum).0.uncertainityBit\ := False;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.34\ := \Unum::AddExactUnums(Unum,Unum).0.num3\ < to_signed(0, 32);
                            \Unum::AddExactUnums(Unum,Unum).0.flag10\ := \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.34\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_132\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_132\.
                            --     * The false branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_133\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_134\.
                            --     * Execution after either branch will continue in the following state: \Unum::AddExactUnums(Unum,Unum).0._State_131\.

                            if (\Unum::AddExactUnums(Unum,Unum).0.flag10\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_132\;
                            else 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_133\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_131\ => 
                        -- State after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_130\.
                        \Unum::AddExactUnums(Unum,Unum).0.num5\ := to_unsigned(0, 16);
                        -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.BitMask::GetMostSignificantOnePosition()
                        \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.bitMask\;
                        \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_135\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_132\ => 
                        -- True branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_130\.
                        \Unum::AddExactUnums(Unum,Unum).0.uncertainityBit\ := True;
                        -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_130\.
                        if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_132\) then 
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_131\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_133\ => 
                        -- False branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_130\.
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::ShiftOutLeastSignificantZeros()
                        \Unum::AddExactUnums(Unum,Unum).0.BitMask::ShiftOutLeastSignificantZeros().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.bitMask\;
                        \Unum::AddExactUnums(Unum,Unum).0.BitMask::ShiftOutLeastSignificantZeros()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_134\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_134\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::ShiftOutLeastSignificantZeros()
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::ShiftOutLeastSignificantZeros()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.BitMask::ShiftOutLeastSignificantZeros()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::ShiftOutLeastSignificantZeros()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.66\ := \Unum::AddExactUnums(Unum,Unum).0.BitMask::ShiftOutLeastSignificantZeros().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.bitMask\ := \Unum::AddExactUnums(Unum,Unum).0.return.66\;
                            -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_130\.
                            if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_134\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_131\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_135\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.BitMask::GetMostSignificantOnePosition()
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.67\ := \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.35\ := \Unum::AddExactUnums(Unum,Unum).0.return.67\ = to_unsigned(0, 16);
                            \Unum::AddExactUnums(Unum,Unum).0.flag11\ := \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.35\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_137\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_137\.
                            --     * The false branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_138\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_139\.
                            --     * Execution after either branch will continue in the following state: \Unum::AddExactUnums(Unum,Unum).0._State_136\.

                            if (\Unum::AddExactUnums(Unum,Unum).0.flag11\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_137\;
                            else 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_138\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_136\ => 
                        -- State after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_135\.
                        -- The last invocation for the target state machine finished in the previous state, so need to start the next one in the next state.
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_140\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_137\ => 
                        -- True branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_135\.
                        \Unum::AddExactUnums(Unum,Unum).0.exponent\ := \Unum::AddExactUnums(Unum,Unum).0.bitMask\;
                        \Unum::AddExactUnums(Unum,Unum).0.exponentSize\ := to_unsigned(0, 8);
                        -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_135\.
                        if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_137\) then 
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_136\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_138\ => 
                        -- False branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_135\.
                        -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.BitMask::GetMostSignificantOnePosition()
                        \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.bitMask\;
                        \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_139\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_139\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.BitMask::GetMostSignificantOnePosition()
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.68\ := \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.36\ := \Unum::AddExactUnums(Unum,Unum).0.return.68\ - to_unsigned(1, 16);
                            \Unum::AddExactUnums(Unum,Unum).0.num5\ := \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.36\;
                            -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_135\.
                            if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_139\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_136\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_140\ => 
                        -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.BitMask::GetMostSignificantOnePosition()
                        \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.exponent\;
                        \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_141\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_141\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.BitMask::GetMostSignificantOnePosition()
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.69\ := \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.37\ := \Unum::AddExactUnums(Unum,Unum).0.return.69\ > to_unsigned(0, 16);
                            \Unum::AddExactUnums(Unum,Unum).0.flag12\ := \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.37\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_143\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_146\.
                            --     * Execution after either branch will continue in the following state: \Unum::AddExactUnums(Unum,Unum).0._State_142\.

                            if (\Unum::AddExactUnums(Unum,Unum).0.flag12\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_143\;
                            else 
                                -- There was no false branch, so going directly to the state after the if-else.
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_142\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_142\ => 
                        -- State after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_141\.
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::IsExact()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsExact().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.left\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsExact()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_149\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_143\ => 
                        -- True branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_141\.
                        -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.BitMask::GetMostSignificantOnePosition()
                        \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.bitMask\;
                        \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_144\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_144\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.BitMask::GetMostSignificantOnePosition()
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.70\ := \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.38\ := \Unum::AddExactUnums(Unum,Unum).0.return.70\ - to_unsigned(1, 16);
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetZero(System.UInt16)
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::SetZero(UInt16).this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.bitMask\;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::SetZero(UInt16).index.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.38\;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::SetZero(UInt16)._Started.0\ <= true;
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_145\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_145\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetZero(System.UInt16)
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::SetZero(UInt16)._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.BitMask::SetZero(UInt16)._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::SetZero(UInt16)._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.71\ := \Unum::AddExactUnums(Unum,Unum).0.BitMask::SetZero(UInt16).return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.bitMask\ := \Unum::AddExactUnums(Unum,Unum).0.return.71\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.39\ := \Unum::AddExactUnums(Unum,Unum).0.num5\ = to_unsigned(0, 16);

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_147\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_147\.
                            --     * The false branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_148\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_148\.
                            --     * Execution after either branch will continue in the following state: \Unum::AddExactUnums(Unum,Unum).0._State_146\.

                            if (\Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.39\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_147\;
                            else 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_148\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_146\ => 
                        -- State after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_145\.
                        -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_141\.
                        if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_146\) then 
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_142\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_147\ => 
                        -- True branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_145\.
                        \Unum::AddExactUnums(Unum,Unum).0.num5\ := to_unsigned(0, 16);
                        -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_145\.
                        if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_147\) then 
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_146\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_148\ => 
                        -- False branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_145\.
                        \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.40\ := \Unum::AddExactUnums(Unum,Unum).0.num5\ - to_unsigned(1, 16);
                        \Unum::AddExactUnums(Unum,Unum).0.num5\ := \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.40\;
                        -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_145\.
                        if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_148\) then 
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_146\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_149\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::IsExact()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::IsExact()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::IsExact()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsExact()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.72\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::IsExact().return.0\;
                            -- The last invocation for the target state machine just finished, so need to start the next one in a later state.
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_150\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_150\ => 
                        -- This state was just added to leave time for the invocation proxy to register that the previous invocation finished.
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_151\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_151\ => 
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.Unum::IsExact()
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsExact().this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.right\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::IsExact()._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_152\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_152\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.Unum::IsExact()
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::IsExact()._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::IsExact()._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsExact()._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.73\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::IsExact().return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.41\ := not(\Unum::AddExactUnums(Unum,Unum).0.return.72\) or not(\Unum::AddExactUnums(Unum,Unum).0.return.73\);
                            \Unum::AddExactUnums(Unum,Unum).0.flag13\ := \Unum::AddExactUnums(Unum,Unum).0.binaryOperationResult.41\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::AddExactUnums(Unum,Unum).0._State_154\ and ends in state \Unum::AddExactUnums(Unum,Unum).0._State_154\.
                            --     * Execution after either branch will continue in the following state: \Unum::AddExactUnums(Unum,Unum).0._State_153\.

                            if (\Unum::AddExactUnums(Unum,Unum).0.flag13\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_154\;
                            else 
                                -- There was no false branch, so going directly to the state after the if-else.
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_153\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::AddExactUnums(Unum,Unum).0._State_153\ => 
                        -- State after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_152\.
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.Unum::SetUnumBits(System.Boolean,Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean,System.Byte,System.UInt16)
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).this.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.unum\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).signBit.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.signBit\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).exponent.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.exponent\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).fraction.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.bitMask\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).uncertainityBit.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.uncertainityBit\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).exponentSize.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.exponentSize\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).fractionSize.parameter.Out.0\ <= \Unum::AddExactUnums(Unum,Unum).0.num5\;
                        \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Started.0\ <= true;
                        \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_155\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_154\ => 
                        -- True branch of the if-else started in state \Unum::AddExactUnums(Unum,Unum).0._State_152\.
                        \Unum::AddExactUnums(Unum,Unum).0.uncertainityBit\ := True;
                        -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_152\.
                        if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_154\) then 
                            \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_153\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddExactUnums(Unum,Unum).0._State_155\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.Unum::SetUnumBits(System.Boolean,Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean,System.Byte,System.UInt16)
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Started.0\ = \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Finished.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Started.0\ <= false;
                            \Unum::AddExactUnums(Unum,Unum).0.return.74\ := \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).return.0\;
                            \Unum::AddExactUnums(Unum,Unum).0.unum\.\UnumBits\ := \Unum::AddExactUnums(Unum,Unum).0.return.74\;
                            \Unum::AddExactUnums(Unum,Unum).0.result\ := \Unum::AddExactUnums(Unum,Unum).0.unum\;
                            -- Going to the state after the if-else which was started in state \Unum::AddExactUnums(Unum,Unum).0._State_36\.
                            if (\Unum::AddExactUnums(Unum,Unum).0._State\ = \Unum::AddExactUnums(Unum,Unum).0._State_155\) then 
                                \Unum::AddExactUnums(Unum,Unum).0._State\ := \Unum::AddExactUnums(Unum,Unum).0._State_37\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentValueToExponentBits(System.Int32,System.Byte).0 state machine start
    \Unum::ExponentValueToExponentBits(Int32,Byte).0._StateMachine\: process (\Clock\) 
        Variable \Unum::ExponentValueToExponentBits(Int32,Byte).0._State\: \Unum::ExponentValueToExponentBits(Int32,Byte).0._States\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_0\;
        Variable \Unum::ExponentValueToExponentBits(Int32,Byte).0.value\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Unum::ExponentValueToExponentBits(Int32,Byte).0.size\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Unum::ExponentValueToExponentBits(Int32,Byte).0.flag\: boolean := false;
        Variable \Unum::ExponentValueToExponentBits(Int32,Byte).0.bitMask\: \Lombiq.Unum.BitMask\;
        Variable \Unum::ExponentValueToExponentBits(Int32,Byte).0.b\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Unum::ExponentValueToExponentBits(Int32,Byte).0.result\: \Lombiq.Unum.BitMask\;
        Variable \Unum::ExponentValueToExponentBits(Int32,Byte).0.bitMask2\: \Lombiq.Unum.BitMask\;
        Variable \Unum::ExponentValueToExponentBits(Int32,Byte).0.b2\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Unum::ExponentValueToExponentBits(Int32,Byte).0.binaryOperationResult.0\: boolean := false;
        Variable \Unum::ExponentValueToExponentBits(Int32,Byte).0.arrayb13ad85d0ff1fab74968cf9635ef50690e8d16091f4b3f34e92839feb21f4e4b\: \unsigned32_Array\(0 to 0) := (others => to_unsigned(0, 32));
        Variable \Unum::ExponentValueToExponentBits(Int32,Byte).0.return.0\: \Lombiq.Unum.BitMask\;
        Variable \Unum::ExponentValueToExponentBits(Int32,Byte).0.array7a549cf35ad1845b7d5eda1814cfb58f101387923beef79cb543eb08d8bec093\: \unsigned32_Array\(0 to 0) := (others => to_unsigned(0, 32));
        Variable \Unum::ExponentValueToExponentBits(Int32,Byte).0.return.1\: \Lombiq.Unum.BitMask\;
        Variable \Unum::ExponentValueToExponentBits(Int32,Byte).0.binaryOperationResult.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Unum::ExponentValueToExponentBits(Int32,Byte).0.return.2\: \Lombiq.Unum.BitMask\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::ExponentValueToExponentBits(Int32,Byte).0._Finished\ <= false;
                \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 32));
                \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\ <= to_unsigned(0, 32);
                \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ <= false;
                \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).right.parameter.Out.0\ <= to_unsigned(0, 32);
                \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ <= false;
                \Unum::ExponentValueToExponentBits(Int32,Byte).0._State\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_0\;
                \Unum::ExponentValueToExponentBits(Int32,Byte).0.value\ := to_signed(0, 32);
                \Unum::ExponentValueToExponentBits(Int32,Byte).0.size\ := to_unsigned(0, 8);
                \Unum::ExponentValueToExponentBits(Int32,Byte).0.flag\ := false;
                \Unum::ExponentValueToExponentBits(Int32,Byte).0.b\ := to_unsigned(0, 8);
                \Unum::ExponentValueToExponentBits(Int32,Byte).0.b2\ := to_unsigned(0, 8);
                \Unum::ExponentValueToExponentBits(Int32,Byte).0.binaryOperationResult.0\ := false;
                \Unum::ExponentValueToExponentBits(Int32,Byte).0.arrayb13ad85d0ff1fab74968cf9635ef50690e8d16091f4b3f34e92839feb21f4e4b\ := (others => to_unsigned(0, 32));
                \Unum::ExponentValueToExponentBits(Int32,Byte).0.array7a549cf35ad1845b7d5eda1814cfb58f101387923beef79cb543eb08d8bec093\ := (others => to_unsigned(0, 32));
                \Unum::ExponentValueToExponentBits(Int32,Byte).0.binaryOperationResult.1\ := to_unsigned(0, 32);
            else 
                case \Unum::ExponentValueToExponentBits(Int32,Byte).0._State\ is 
                    when \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::ExponentValueToExponentBits(Int32,Byte).0._Started\ = true) then 
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0._State\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::ExponentValueToExponentBits(Int32,Byte).0._Started\ = true) then 
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0._Finished\ <= true;
                        else 
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0._Finished\ <= false;
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0._State\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_2\ => 
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.value\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0.value.parameter.In\;
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.size\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0.size.parameter.In\;
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.binaryOperationResult.0\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0.value\ > to_signed(0, 32);
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.flag\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0.binaryOperationResult.0\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_4\ and ends in state \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_6\.
                        --     * The false branch starts in state \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_7\ and ends in state \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_10\.
                        --     * Execution after either branch will continue in the following state: \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_3\.

                        if (\Unum::ExponentValueToExponentBits(Int32,Byte).0.flag\) then 
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0._State\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_4\;
                        else 
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0._State\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_3\ => 
                        -- State after the if-else which was started in state \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_2\.
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.return\ <= \Unum::ExponentValueToExponentBits(Int32,Byte).0.result\;
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0._State\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_4\ => 
                        -- True branch of the if-else started in state \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_2\.
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.arrayb13ad85d0ff1fab74968cf9635ef50690e8d16091f4b3f34e92839feb21f4e4b\ := (others => to_unsigned(0, 32));
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.arrayb13ad85d0ff1fab74968cf9635ef50690e8d16091f4b3f34e92839feb21f4e4b\(to_integer(to_signed(0, 32))) := unsigned(\Unum::ExponentValueToExponentBits(Int32,Byte).0.value\);
                        -- Initializing record fields to their defaults.
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.bitMask\.\IsNull\ := false;
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.bitMask\.\Size\ := to_unsigned(0, 16);
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.bitMask\.\SegmentCount\ := to_unsigned(0, 16);
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.bitMask\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\ <= \Unum::ExponentValueToExponentBits(Int32,Byte).0.bitMask\;
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\(0 to 0) <= \Unum::ExponentValueToExponentBits(Int32,Byte).0.arrayb13ad85d0ff1fab74968cf9635ef50690e8d16091f4b3f34e92839feb21f4e4b\;
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= resize(\Unum::ExponentValueToExponentBits(Int32,Byte).0.size\, 16);
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= true;
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0._State\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_5\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        if (\Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\) then 
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.bitMask\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\;
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.arrayb13ad85d0ff1fab74968cf9635ef50690e8d16091f4b3f34e92839feb21f4e4b\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\(0 to 0);
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.b\ := to_unsigned(1, 8);
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,System.UInt32)
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32).left.parameter.Out.0\ <= \Unum::ExponentValueToExponentBits(Int32,Byte).0.bitMask\;
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\ <= to_unsigned(0, 32);
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ <= true;
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0._State\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_6\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,System.UInt32)
                        if (\Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ = \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\) then 
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ <= false;
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.return.0\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32).return.0\;
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.bitMask\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0.return.0\;
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.result\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0.bitMask\;
                            -- Going to the state after the if-else which was started in state \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_2\.
                            if (\Unum::ExponentValueToExponentBits(Int32,Byte).0._State\ = \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_6\) then 
                                \Unum::ExponentValueToExponentBits(Int32,Byte).0._State\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_3\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_7\ => 
                        -- False branch of the if-else started in state \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_2\.
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.array7a549cf35ad1845b7d5eda1814cfb58f101387923beef79cb543eb08d8bec093\ := (others => to_unsigned(0, 32));
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.array7a549cf35ad1845b7d5eda1814cfb58f101387923beef79cb543eb08d8bec093\(to_integer(to_signed(0, 32))) := unsigned(signed(0 - unsigned(\Unum::ExponentValueToExponentBits(Int32,Byte).0.value\)));
                        -- Initializing record fields to their defaults.
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.bitMask2\.\IsNull\ := false;
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.bitMask2\.\Size\ := to_unsigned(0, 16);
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.bitMask2\.\SegmentCount\ := to_unsigned(0, 16);
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.bitMask2\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\ <= \Unum::ExponentValueToExponentBits(Int32,Byte).0.bitMask2\;
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\(0 to 0) <= \Unum::ExponentValueToExponentBits(Int32,Byte).0.array7a549cf35ad1845b7d5eda1814cfb58f101387923beef79cb543eb08d8bec093\;
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\ <= resize(\Unum::ExponentValueToExponentBits(Int32,Byte).0.size\, 16);
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= true;
                        \Unum::ExponentValueToExponentBits(Int32,Byte).0._State\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_8\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_8\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16)
                        if (\Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\) then 
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ <= false;
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.bitMask2\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\;
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.array7a549cf35ad1845b7d5eda1814cfb58f101387923beef79cb543eb08d8bec093\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\(0 to 0);
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.b2\ := to_unsigned(1, 8);
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,System.UInt32)
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32).left.parameter.Out.0\ <= \Unum::ExponentValueToExponentBits(Int32,Byte).0.bitMask2\;
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\ <= to_unsigned(0, 32);
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ <= true;
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0._State\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_9\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_9\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,System.UInt32)
                        if (\Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ = \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\) then 
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ <= false;
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.return.1\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32).return.0\;
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.bitMask2\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0.return.1\;
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.binaryOperationResult.1\ := resize(unsigned(to_signed(-2, 32) * \Unum::ExponentValueToExponentBits(Int32,Byte).0.value\), 32);
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,System.UInt32)
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).left.parameter.Out.0\ <= \Unum::ExponentValueToExponentBits(Int32,Byte).0.bitMask2\;
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).right.parameter.Out.0\ <= (\Unum::ExponentValueToExponentBits(Int32,Byte).0.binaryOperationResult.1\);
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ <= true;
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0._State\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_10\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_10\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,System.UInt32)
                        if (\Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ = \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\) then 
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ <= false;
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.return.2\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).return.0\;
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.bitMask2\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0.return.2\;
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.result\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0.bitMask2\;
                            -- Going to the state after the if-else which was started in state \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_2\.
                            if (\Unum::ExponentValueToExponentBits(Int32,Byte).0._State\ = \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_10\) then 
                                \Unum::ExponentValueToExponentBits(Int32,Byte).0._State\ := \Unum::ExponentValueToExponentBits(Int32,Byte).0._State_3\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentValueToExponentBits(System.Int32,System.Byte).0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::AddAlignedFractions(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean).0 state machine start
    \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._StateMachine\: process (\Clock\) 
        Variable \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\: \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._States\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_0\;
        Variable \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.left\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.right\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.signBitsMatch\: boolean := false;
        Variable \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.result\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.return.0\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.return.1\: boolean := false;
        Variable \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.return.2\: \Lombiq.Unum.BitMask\;
        Variable \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.return.3\: \Lombiq.Unum.BitMask\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._Finished\ <= false;
                \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\ <= false;
                \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= false;
                \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= false;
                \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_GreaterThan(BitMask,BitMask)._Started.0\ <= false;
                \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ <= false;
                \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_0\;
                \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.signBitsMatch\ := false;
                \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.return.1\ := false;
            else 
                case \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\ is 
                    when \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._Started\ = true) then 
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._Started\ = true) then 
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._Finished\ <= true;
                        else 
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._Finished\ <= false;
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_2\ => 
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.left\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.left.parameter.In\;
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.right\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.right.parameter.In\;
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.signBitsMatch\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.signBitsMatch.parameter.In\;
                        -- Initializing record fields to their defaults.
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.result\.\IsNull\ := false;
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.result\.\Size\ := to_unsigned(0, 16);
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.result\.\SegmentCount\ := to_unsigned(0, 16);
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.result\.\Segments\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\ <= \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.result\;
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\ <= \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.left\.\Size\;
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\ <= False;
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= true;
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                        if (\Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ = \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\) then 
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= false;
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.result\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_5\ and ends in state \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_6\.
                            --     * The false branch starts in state \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_7\ and ends in state \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_9\.
                            --     * Execution after either branch will continue in the following state: \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_4\.

                            if (\Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.signBitsMatch\) then 
                                \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_5\;
                            else 
                                \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_7\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_4\ => 
                        -- State after the if-else which was started in state \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_3\.
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.return\ <= \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.result\;
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_5\ => 
                        -- True branch of the if-else started in state \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_3\.
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Addition(BitMask,BitMask).left.parameter.Out.0\ <= \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.left\;
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Addition(BitMask,BitMask).right.parameter.Out.0\ <= \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.right\;
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= true;
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_6\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_6\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ = \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\) then 
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= false;
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.return.0\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Addition(BitMask,BitMask).return.0\;
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.result\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.return.0\;
                            -- Going to the state after the if-else which was started in state \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_3\.
                            if (\Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\ = \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_6\) then 
                                \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_4\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_7\ => 
                        -- False branch of the if-else started in state \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_3\.
                        -- Starting state machine invocation for the following method: System.Boolean Lombiq.Unum.BitMask::op_GreaterThan(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_GreaterThan(BitMask,BitMask).left.parameter.Out.0\ <= \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.left\;
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_GreaterThan(BitMask,BitMask).right.parameter.Out.0\ <= \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.right\;
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_GreaterThan(BitMask,BitMask)._Started.0\ <= true;
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_8\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_8\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Lombiq.Unum.BitMask::op_GreaterThan(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_GreaterThan(BitMask,BitMask)._Started.0\ = \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_GreaterThan(BitMask,BitMask)._Finished.0\) then 
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_GreaterThan(BitMask,BitMask)._Started.0\ <= false;
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.return.1\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_GreaterThan(BitMask,BitMask).return.0\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_10\ and ends in state \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_11\.
                            --     * The false branch starts in state \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_12\ and ends in state \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_14\.
                            --     * Execution after either branch will continue in the following state: \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_9\.

                            if (\Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.return.1\) then 
                                \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_10\;
                            else 
                                \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_12\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_9\ => 
                        -- State after the if-else which was started in state \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_8\.
                        -- Going to the state after the if-else which was started in state \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_3\.
                        if (\Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\ = \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_9\) then 
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_10\ => 
                        -- True branch of the if-else started in state \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_8\.
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask).left.parameter.Out.0\ <= \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.left\;
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask).right.parameter.Out.0\ <= \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.right\;
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ <= true;
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_11\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_11\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ = \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask)._Finished.0\) then 
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ <= false;
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.return.2\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask).return.0\;
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.result\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.return.2\;
                            -- Going to the state after the if-else which was started in state \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_8\.
                            if (\Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\ = \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_11\) then 
                                \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_9\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_12\ => 
                        -- False branch of the if-else started in state \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_8\.
                        -- The last invocation for the target state machine finished in the previous state, so need to start the next one in the next state.
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_13\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_13\ => 
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask).left.parameter.Out.0\ <= \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.right\;
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask).right.parameter.Out.0\ <= \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.left\;
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ <= true;
                        \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_14\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_14\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ = \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask)._Finished.0\) then 
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ <= false;
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.return.3\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask).return.0\;
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.result\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.return.3\;
                            -- Going to the state after the if-else which was started in state \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_8\.
                            if (\Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\ = \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_14\) then 
                                \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State\ := \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._State_9\;
                            end if;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::AddAlignedFractions(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean).0 state machine end


    -- Lombiq.Unum.Unum Lombiq.Unum.Unum::op_Addition(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0 state machine start
    \Unum::op_Addition(Unum,Unum).0._StateMachine\: process (\Clock\) 
        Variable \Unum::op_Addition(Unum,Unum).0._State\: \Unum::op_Addition(Unum,Unum).0._States\ := \Unum::op_Addition(Unum,Unum).0._State_0\;
        Variable \Unum::op_Addition(Unum,Unum).0.left\: \Lombiq.Unum.Unum\;
        Variable \Unum::op_Addition(Unum,Unum).0.right\: \Lombiq.Unum.Unum\;
        Variable \Unum::op_Addition(Unum,Unum).0.return.0\: \Lombiq.Unum.Unum\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::op_Addition(Unum,Unum).0._Finished\ <= false;
                \Unum::op_Addition(Unum,Unum).0.Unum::AddExactUnums(Unum,Unum)._Started.0\ <= false;
                \Unum::op_Addition(Unum,Unum).0._State\ := \Unum::op_Addition(Unum,Unum).0._State_0\;
            else 
                case \Unum::op_Addition(Unum,Unum).0._State\ is 
                    when \Unum::op_Addition(Unum,Unum).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::op_Addition(Unum,Unum).0._Started\ = true) then 
                            \Unum::op_Addition(Unum,Unum).0._State\ := \Unum::op_Addition(Unum,Unum).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::op_Addition(Unum,Unum).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::op_Addition(Unum,Unum).0._Started\ = true) then 
                            \Unum::op_Addition(Unum,Unum).0._Finished\ <= true;
                        else 
                            \Unum::op_Addition(Unum,Unum).0._Finished\ <= false;
                            \Unum::op_Addition(Unum,Unum).0._State\ := \Unum::op_Addition(Unum,Unum).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::op_Addition(Unum,Unum).0._State_2\ => 
                        \Unum::op_Addition(Unum,Unum).0.left\ := \Unum::op_Addition(Unum,Unum).0.left.parameter.In\;
                        \Unum::op_Addition(Unum,Unum).0.right\ := \Unum::op_Addition(Unum,Unum).0.right.parameter.In\;
                        -- Starting state machine invocation for the following method: Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum)
                        \Unum::op_Addition(Unum,Unum).0.Unum::AddExactUnums(Unum,Unum).left.parameter.Out.0\ <= \Unum::op_Addition(Unum,Unum).0.left\;
                        \Unum::op_Addition(Unum,Unum).0.Unum::AddExactUnums(Unum,Unum).right.parameter.Out.0\ <= \Unum::op_Addition(Unum,Unum).0.right\;
                        \Unum::op_Addition(Unum,Unum).0.Unum::AddExactUnums(Unum,Unum)._Started.0\ <= true;
                        \Unum::op_Addition(Unum,Unum).0._State\ := \Unum::op_Addition(Unum,Unum).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::op_Addition(Unum,Unum).0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum)
                        if (\Unum::op_Addition(Unum,Unum).0.Unum::AddExactUnums(Unum,Unum)._Started.0\ = \Unum::op_Addition(Unum,Unum).0.Unum::AddExactUnums(Unum,Unum)._Finished.0\) then 
                            \Unum::op_Addition(Unum,Unum).0.Unum::AddExactUnums(Unum,Unum)._Started.0\ <= false;
                            \Unum::op_Addition(Unum,Unum).0.return.0\ := \Unum::op_Addition(Unum,Unum).0.Unum::AddExactUnums(Unum,Unum).return.0\;
                            \Unum::op_Addition(Unum,Unum).0.return\ <= \Unum::op_Addition(Unum,Unum).0.return.0\;
                            \Unum::op_Addition(Unum,Unum).0._State\ := \Unum::op_Addition(Unum,Unum).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.Unum Lombiq.Unum.Unum::op_Addition(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0 state machine end


    -- System.UInt16 Lombiq.Unum.Unum::get_FractionSizeMax().0 state machine start
    \Unum::get_FractionSizeMax().0._StateMachine\: process (\Clock\) 
        Variable \Unum::get_FractionSizeMax().0._State\: \Unum::get_FractionSizeMax().0._States\ := \Unum::get_FractionSizeMax().0._State_0\;
        Variable \Unum::get_FractionSizeMax().0.this\: \Lombiq.Unum.Unum\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::get_FractionSizeMax().0._Finished\ <= false;
                \Unum::get_FractionSizeMax().0.return\ <= to_unsigned(0, 16);
                \Unum::get_FractionSizeMax().0._State\ := \Unum::get_FractionSizeMax().0._State_0\;
            else 
                case \Unum::get_FractionSizeMax().0._State\ is 
                    when \Unum::get_FractionSizeMax().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::get_FractionSizeMax().0._Started\ = true) then 
                            \Unum::get_FractionSizeMax().0._State\ := \Unum::get_FractionSizeMax().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::get_FractionSizeMax().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::get_FractionSizeMax().0._Started\ = true) then 
                            \Unum::get_FractionSizeMax().0._Finished\ <= true;
                        else 
                            \Unum::get_FractionSizeMax().0._Finished\ <= false;
                            \Unum::get_FractionSizeMax().0._State\ := \Unum::get_FractionSizeMax().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::get_FractionSizeMax().0._State_2\ => 
                        \Unum::get_FractionSizeMax().0.this\ := \Unum::get_FractionSizeMax().0.this.parameter.In\;
                        \Unum::get_FractionSizeMax().0.return\ <= \Unum::get_FractionSizeMax().0.this\.\_environment\.\FractionSizeMax\;
                        \Unum::get_FractionSizeMax().0._State\ := \Unum::get_FractionSizeMax().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.UInt16 Lombiq.Unum.Unum::get_FractionSizeMax().0 state machine end


    -- System.UInt16 Lombiq.Unum.Unum::get_Size().0 state machine start
    \Unum::get_Size().0._StateMachine\: process (\Clock\) 
        Variable \Unum::get_Size().0._State\: \Unum::get_Size().0._States\ := \Unum::get_Size().0._State_0\;
        Variable \Unum::get_Size().0.this\: \Lombiq.Unum.Unum\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::get_Size().0._Finished\ <= false;
                \Unum::get_Size().0.return\ <= to_unsigned(0, 16);
                \Unum::get_Size().0._State\ := \Unum::get_Size().0._State_0\;
            else 
                case \Unum::get_Size().0._State\ is 
                    when \Unum::get_Size().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::get_Size().0._Started\ = true) then 
                            \Unum::get_Size().0._State\ := \Unum::get_Size().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::get_Size().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::get_Size().0._Started\ = true) then 
                            \Unum::get_Size().0._Finished\ <= true;
                        else 
                            \Unum::get_Size().0._Finished\ <= false;
                            \Unum::get_Size().0._State\ := \Unum::get_Size().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::get_Size().0._State_2\ => 
                        \Unum::get_Size().0.this\ := \Unum::get_Size().0.this.parameter.In\;
                        \Unum::get_Size().0.return\ <= \Unum::get_Size().0.this\.\_environment\.\Size\;
                        \Unum::get_Size().0._State\ := \Unum::get_Size().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.UInt16 Lombiq.Unum.Unum::get_Size().0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_UncertaintyBitMask().0 state machine start
    \Unum::get_UncertaintyBitMask().0._StateMachine\: process (\Clock\) 
        Variable \Unum::get_UncertaintyBitMask().0._State\: \Unum::get_UncertaintyBitMask().0._States\ := \Unum::get_UncertaintyBitMask().0._State_0\;
        Variable \Unum::get_UncertaintyBitMask().0.this\: \Lombiq.Unum.Unum\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::get_UncertaintyBitMask().0._Finished\ <= false;
                \Unum::get_UncertaintyBitMask().0._State\ := \Unum::get_UncertaintyBitMask().0._State_0\;
            else 
                case \Unum::get_UncertaintyBitMask().0._State\ is 
                    when \Unum::get_UncertaintyBitMask().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::get_UncertaintyBitMask().0._Started\ = true) then 
                            \Unum::get_UncertaintyBitMask().0._State\ := \Unum::get_UncertaintyBitMask().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::get_UncertaintyBitMask().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::get_UncertaintyBitMask().0._Started\ = true) then 
                            \Unum::get_UncertaintyBitMask().0._Finished\ <= true;
                        else 
                            \Unum::get_UncertaintyBitMask().0._Finished\ <= false;
                            \Unum::get_UncertaintyBitMask().0._State\ := \Unum::get_UncertaintyBitMask().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::get_UncertaintyBitMask().0._State_2\ => 
                        \Unum::get_UncertaintyBitMask().0.this\ := \Unum::get_UncertaintyBitMask().0.this.parameter.In\;
                        \Unum::get_UncertaintyBitMask().0.return\ <= \Unum::get_UncertaintyBitMask().0.this\.\_environment\.\UncertaintyBitMask\;
                        \Unum::get_UncertaintyBitMask().0._State\ := \Unum::get_UncertaintyBitMask().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_UncertaintyBitMask().0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_ExponentSizeMask().0 state machine start
    \Unum::get_ExponentSizeMask().0._StateMachine\: process (\Clock\) 
        Variable \Unum::get_ExponentSizeMask().0._State\: \Unum::get_ExponentSizeMask().0._States\ := \Unum::get_ExponentSizeMask().0._State_0\;
        Variable \Unum::get_ExponentSizeMask().0.this\: \Lombiq.Unum.Unum\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::get_ExponentSizeMask().0._Finished\ <= false;
                \Unum::get_ExponentSizeMask().0._State\ := \Unum::get_ExponentSizeMask().0._State_0\;
            else 
                case \Unum::get_ExponentSizeMask().0._State\ is 
                    when \Unum::get_ExponentSizeMask().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::get_ExponentSizeMask().0._Started\ = true) then 
                            \Unum::get_ExponentSizeMask().0._State\ := \Unum::get_ExponentSizeMask().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::get_ExponentSizeMask().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::get_ExponentSizeMask().0._Started\ = true) then 
                            \Unum::get_ExponentSizeMask().0._Finished\ <= true;
                        else 
                            \Unum::get_ExponentSizeMask().0._Finished\ <= false;
                            \Unum::get_ExponentSizeMask().0._State\ := \Unum::get_ExponentSizeMask().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::get_ExponentSizeMask().0._State_2\ => 
                        \Unum::get_ExponentSizeMask().0.this\ := \Unum::get_ExponentSizeMask().0.this.parameter.In\;
                        \Unum::get_ExponentSizeMask().0.return\ <= \Unum::get_ExponentSizeMask().0.this\.\_environment\.\ExponentSizeMask\;
                        \Unum::get_ExponentSizeMask().0._State\ := \Unum::get_ExponentSizeMask().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_ExponentSizeMask().0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_FractionSizeMask().0 state machine start
    \Unum::get_FractionSizeMask().0._StateMachine\: process (\Clock\) 
        Variable \Unum::get_FractionSizeMask().0._State\: \Unum::get_FractionSizeMask().0._States\ := \Unum::get_FractionSizeMask().0._State_0\;
        Variable \Unum::get_FractionSizeMask().0.this\: \Lombiq.Unum.Unum\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::get_FractionSizeMask().0._Finished\ <= false;
                \Unum::get_FractionSizeMask().0._State\ := \Unum::get_FractionSizeMask().0._State_0\;
            else 
                case \Unum::get_FractionSizeMask().0._State\ is 
                    when \Unum::get_FractionSizeMask().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::get_FractionSizeMask().0._Started\ = true) then 
                            \Unum::get_FractionSizeMask().0._State\ := \Unum::get_FractionSizeMask().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::get_FractionSizeMask().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::get_FractionSizeMask().0._Started\ = true) then 
                            \Unum::get_FractionSizeMask().0._Finished\ <= true;
                        else 
                            \Unum::get_FractionSizeMask().0._Finished\ <= false;
                            \Unum::get_FractionSizeMask().0._State\ := \Unum::get_FractionSizeMask().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::get_FractionSizeMask().0._State_2\ => 
                        \Unum::get_FractionSizeMask().0.this\ := \Unum::get_FractionSizeMask().0.this.parameter.In\;
                        \Unum::get_FractionSizeMask().0.return\ <= \Unum::get_FractionSizeMask().0.this\.\_environment\.\FractionSizeMask\;
                        \Unum::get_FractionSizeMask().0._State\ := \Unum::get_FractionSizeMask().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_FractionSizeMask().0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_SignBitMask().0 state machine start
    \Unum::get_SignBitMask().0._StateMachine\: process (\Clock\) 
        Variable \Unum::get_SignBitMask().0._State\: \Unum::get_SignBitMask().0._States\ := \Unum::get_SignBitMask().0._State_0\;
        Variable \Unum::get_SignBitMask().0.this\: \Lombiq.Unum.Unum\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::get_SignBitMask().0._Finished\ <= false;
                \Unum::get_SignBitMask().0._State\ := \Unum::get_SignBitMask().0._State_0\;
            else 
                case \Unum::get_SignBitMask().0._State\ is 
                    when \Unum::get_SignBitMask().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::get_SignBitMask().0._Started\ = true) then 
                            \Unum::get_SignBitMask().0._State\ := \Unum::get_SignBitMask().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::get_SignBitMask().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::get_SignBitMask().0._Started\ = true) then 
                            \Unum::get_SignBitMask().0._Finished\ <= true;
                        else 
                            \Unum::get_SignBitMask().0._Finished\ <= false;
                            \Unum::get_SignBitMask().0._State\ := \Unum::get_SignBitMask().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::get_SignBitMask().0._State_2\ => 
                        \Unum::get_SignBitMask().0.this\ := \Unum::get_SignBitMask().0.this.parameter.In\;
                        \Unum::get_SignBitMask().0.return\ <= \Unum::get_SignBitMask().0.this\.\_environment\.\SignBitMask\;
                        \Unum::get_SignBitMask().0._State\ := \Unum::get_SignBitMask().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_SignBitMask().0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_PositiveInfinity().0 state machine start
    \Unum::get_PositiveInfinity().0._StateMachine\: process (\Clock\) 
        Variable \Unum::get_PositiveInfinity().0._State\: \Unum::get_PositiveInfinity().0._States\ := \Unum::get_PositiveInfinity().0._State_0\;
        Variable \Unum::get_PositiveInfinity().0.this\: \Lombiq.Unum.Unum\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::get_PositiveInfinity().0._Finished\ <= false;
                \Unum::get_PositiveInfinity().0._State\ := \Unum::get_PositiveInfinity().0._State_0\;
            else 
                case \Unum::get_PositiveInfinity().0._State\ is 
                    when \Unum::get_PositiveInfinity().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::get_PositiveInfinity().0._Started\ = true) then 
                            \Unum::get_PositiveInfinity().0._State\ := \Unum::get_PositiveInfinity().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::get_PositiveInfinity().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::get_PositiveInfinity().0._Started\ = true) then 
                            \Unum::get_PositiveInfinity().0._Finished\ <= true;
                        else 
                            \Unum::get_PositiveInfinity().0._Finished\ <= false;
                            \Unum::get_PositiveInfinity().0._State\ := \Unum::get_PositiveInfinity().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::get_PositiveInfinity().0._State_2\ => 
                        \Unum::get_PositiveInfinity().0.this\ := \Unum::get_PositiveInfinity().0.this.parameter.In\;
                        \Unum::get_PositiveInfinity().0.return\ <= \Unum::get_PositiveInfinity().0.this\.\_environment\.\PositiveInfinity\;
                        \Unum::get_PositiveInfinity().0._State\ := \Unum::get_PositiveInfinity().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_PositiveInfinity().0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_NegativeInfinity().0 state machine start
    \Unum::get_NegativeInfinity().0._StateMachine\: process (\Clock\) 
        Variable \Unum::get_NegativeInfinity().0._State\: \Unum::get_NegativeInfinity().0._States\ := \Unum::get_NegativeInfinity().0._State_0\;
        Variable \Unum::get_NegativeInfinity().0.this\: \Lombiq.Unum.Unum\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::get_NegativeInfinity().0._Finished\ <= false;
                \Unum::get_NegativeInfinity().0._State\ := \Unum::get_NegativeInfinity().0._State_0\;
            else 
                case \Unum::get_NegativeInfinity().0._State\ is 
                    when \Unum::get_NegativeInfinity().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::get_NegativeInfinity().0._Started\ = true) then 
                            \Unum::get_NegativeInfinity().0._State\ := \Unum::get_NegativeInfinity().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::get_NegativeInfinity().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::get_NegativeInfinity().0._Started\ = true) then 
                            \Unum::get_NegativeInfinity().0._Finished\ <= true;
                        else 
                            \Unum::get_NegativeInfinity().0._Finished\ <= false;
                            \Unum::get_NegativeInfinity().0._State\ := \Unum::get_NegativeInfinity().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::get_NegativeInfinity().0._State_2\ => 
                        \Unum::get_NegativeInfinity().0.this\ := \Unum::get_NegativeInfinity().0.this.parameter.In\;
                        \Unum::get_NegativeInfinity().0.return\ <= \Unum::get_NegativeInfinity().0.this\.\_environment\.\NegativeInfinity\;
                        \Unum::get_NegativeInfinity().0._State\ := \Unum::get_NegativeInfinity().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_NegativeInfinity().0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_QuietNotANumber().0 state machine start
    \Unum::get_QuietNotANumber().0._StateMachine\: process (\Clock\) 
        Variable \Unum::get_QuietNotANumber().0._State\: \Unum::get_QuietNotANumber().0._States\ := \Unum::get_QuietNotANumber().0._State_0\;
        Variable \Unum::get_QuietNotANumber().0.this\: \Lombiq.Unum.Unum\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::get_QuietNotANumber().0._Finished\ <= false;
                \Unum::get_QuietNotANumber().0._State\ := \Unum::get_QuietNotANumber().0._State_0\;
            else 
                case \Unum::get_QuietNotANumber().0._State\ is 
                    when \Unum::get_QuietNotANumber().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::get_QuietNotANumber().0._Started\ = true) then 
                            \Unum::get_QuietNotANumber().0._State\ := \Unum::get_QuietNotANumber().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::get_QuietNotANumber().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::get_QuietNotANumber().0._Started\ = true) then 
                            \Unum::get_QuietNotANumber().0._Finished\ <= true;
                        else 
                            \Unum::get_QuietNotANumber().0._Finished\ <= false;
                            \Unum::get_QuietNotANumber().0._State\ := \Unum::get_QuietNotANumber().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::get_QuietNotANumber().0._State_2\ => 
                        \Unum::get_QuietNotANumber().0.this\ := \Unum::get_QuietNotANumber().0.this.parameter.In\;
                        \Unum::get_QuietNotANumber().0.return\ <= \Unum::get_QuietNotANumber().0.this\.\_environment\.\QuietNotANumber\;
                        \Unum::get_QuietNotANumber().0._State\ := \Unum::get_QuietNotANumber().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_QuietNotANumber().0 state machine end


    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_SignalingNotANumber().0 state machine start
    \Unum::get_SignalingNotANumber().0._StateMachine\: process (\Clock\) 
        Variable \Unum::get_SignalingNotANumber().0._State\: \Unum::get_SignalingNotANumber().0._States\ := \Unum::get_SignalingNotANumber().0._State_0\;
        Variable \Unum::get_SignalingNotANumber().0.this\: \Lombiq.Unum.Unum\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Unum::get_SignalingNotANumber().0._Finished\ <= false;
                \Unum::get_SignalingNotANumber().0._State\ := \Unum::get_SignalingNotANumber().0._State_0\;
            else 
                case \Unum::get_SignalingNotANumber().0._State\ is 
                    when \Unum::get_SignalingNotANumber().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\Unum::get_SignalingNotANumber().0._Started\ = true) then 
                            \Unum::get_SignalingNotANumber().0._State\ := \Unum::get_SignalingNotANumber().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::get_SignalingNotANumber().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\Unum::get_SignalingNotANumber().0._Started\ = true) then 
                            \Unum::get_SignalingNotANumber().0._Finished\ <= true;
                        else 
                            \Unum::get_SignalingNotANumber().0._Finished\ <= false;
                            \Unum::get_SignalingNotANumber().0._State\ := \Unum::get_SignalingNotANumber().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \Unum::get_SignalingNotANumber().0._State_2\ => 
                        \Unum::get_SignalingNotANumber().0.this\ := \Unum::get_SignalingNotANumber().0.this.parameter.In\;
                        \Unum::get_SignalingNotANumber().0.return\ <= \Unum::get_SignalingNotANumber().0.this\.\_environment\.\SignalingNotANumber\;
                        \Unum::get_SignalingNotANumber().0._State\ := \Unum::get_SignalingNotANumber().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_SignalingNotANumber().0 state machine end


    -- System.UInt16 Lombiq.Unum.UnumHelper::SegmentSizeSizeToSegmentSize(System.Byte).0 state machine start
    \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._StateMachine\: process (\Clock\) 
        Variable \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._State\: \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._States\ := \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._State_0\;
        Variable \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0.segmentSizeSize\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0.binaryOperationResult.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._Finished\ <= false;
                \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0.return\ <= to_unsigned(0, 16);
                \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._State\ := \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._State_0\;
                \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0.segmentSizeSize\ := to_unsigned(0, 8);
                \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0.binaryOperationResult.0\ := to_unsigned(0, 16);
            else 
                case \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._State\ is 
                    when \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._Started\ = true) then 
                            \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._State\ := \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._Started\ = true) then 
                            \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._Finished\ <= true;
                        else 
                            \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._Finished\ <= false;
                            \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._State\ := \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._State_2\ => 
                        \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0.segmentSizeSize\ := \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0.segmentSizeSize.parameter.In\;
                        \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0.binaryOperationResult.0\ := resize(unsigned(shift_left(to_signed(1, 32), to_integer(resize(signed(\UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0.segmentSizeSize\), 32)))), 16);
                        \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0.return\ <= (\UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0.binaryOperationResult.0\);
                        \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._State\ := \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.UInt16 Lombiq.Unum.UnumHelper::SegmentSizeSizeToSegmentSize(System.Byte).0 state machine end


    -- System.Void Lombiq.Unum.UnumEnvironment::.ctor(System.Byte,System.Byte).0 state machine start
    \UnumEnvironment::.ctor(Byte,Byte).0._StateMachine\: process (\Clock\) 
        Variable \UnumEnvironment::.ctor(Byte,Byte).0._State\: \UnumEnvironment::.ctor(Byte,Byte).0._States\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_0\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.this\: \Lombiq.Unum.UnumEnvironment\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.exponentSizeSize\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.fractionSizeSize\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.return.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.return.1\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.1\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.2\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.objecta4c70e00f2ec2975ffd03b87442e75fb219dd43f089d457c217e1f67cffbf4a0\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.return.2\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.object1af8c7e1413e2da44291e3b4786150cb23fed68c0d70afe08a2e21d86ea1dbf3\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.return.3\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.return.4\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.return.5\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.return.6\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.return.7\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.return.8\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.object7f34fefc400743c5659b915282ee58959b74703089d82e84e8d6c948e4b443d7\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.3\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.return.9\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.objecte438b2d1e01c6422c441d4244fd563f19ddf9cd04a02503bb4f07fbb1fcf4864\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.return.10\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.object479fe084fa4366b617a7eeccf1cdebf1ed267e764cb62ef8fe9d94f131cbeab7\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.4\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.return.11\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.return.12\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.return.13\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.objectf4f045d4d2f66a18d2b9627940ae5ecef55676a7cd16373be4c2abd2bc60efc2\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.5\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.return.14\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.return.15\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.return.16\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.return.17\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.return.18\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.6\: signed(31 downto 0) := to_signed(0, 32);
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.7\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.return.19\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.return.20\: \Lombiq.Unum.BitMask\;
        Variable \UnumEnvironment::.ctor(Byte,Byte).0.return.21\: \Lombiq.Unum.BitMask\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \UnumEnvironment::.ctor(Byte,Byte).0._Finished\ <= false;
                \UnumEnvironment::.ctor(Byte,Byte).0.UnumHelper::SegmentSizeSizeToSegmentSize(Byte).segmentSizeSize.parameter.Out.0\ <= to_unsigned(0, 8);
                \UnumEnvironment::.ctor(Byte,Byte).0.UnumHelper::SegmentSizeSizeToSegmentSize(Byte)._Started.0\ <= false;
                \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\ <= false;
                \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= false;
                \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).index.parameter.Out.0\ <= to_unsigned(0, 16);
                \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Started.0\ <= false;
                \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).right.parameter.Out.0\ <= to_unsigned(0, 32);
                \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ <= false;
                \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ <= false;
                \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_BitwiseOr(BitMask,BitMask)._Started.0\ <= false;
                \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= false;
                \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\ <= to_unsigned(0, 32);
                \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ <= false;
                \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_0\;
                \UnumEnvironment::.ctor(Byte,Byte).0.exponentSizeSize\ := to_unsigned(0, 8);
                \UnumEnvironment::.ctor(Byte,Byte).0.fractionSizeSize\ := to_unsigned(0, 8);
                \UnumEnvironment::.ctor(Byte,Byte).0.return.0\ := to_unsigned(0, 16);
                \UnumEnvironment::.ctor(Byte,Byte).0.return.1\ := to_unsigned(0, 16);
                \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.0\ := to_unsigned(0, 16);
                \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.1\ := to_unsigned(0, 16);
                \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.2\ := to_unsigned(0, 16);
                \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.3\ := to_unsigned(0, 16);
                \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.4\ := to_unsigned(0, 16);
                \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.5\ := to_unsigned(0, 16);
                \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.6\ := to_signed(0, 32);
                \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.7\ := to_unsigned(0, 32);
            else 
                case \UnumEnvironment::.ctor(Byte,Byte).0._State\ is 
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\UnumEnvironment::.ctor(Byte,Byte).0._Started\ = true) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\UnumEnvironment::.ctor(Byte,Byte).0._Started\ = true) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0._Finished\ <= true;
                        else 
                            \UnumEnvironment::.ctor(Byte,Byte).0._Finished\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \UnumEnvironment::.ctor(Byte,Byte).0.this.parameter.Out\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_2\ => 
                        \UnumEnvironment::.ctor(Byte,Byte).0.this\ := \UnumEnvironment::.ctor(Byte,Byte).0.this.parameter.In\;
                        \UnumEnvironment::.ctor(Byte,Byte).0.exponentSizeSize\ := \UnumEnvironment::.ctor(Byte,Byte).0.exponentSizeSize.parameter.In\;
                        \UnumEnvironment::.ctor(Byte,Byte).0.fractionSizeSize\ := \UnumEnvironment::.ctor(Byte,Byte).0.fractionSizeSize.parameter.In\;
                        \UnumEnvironment::.ctor(Byte,Byte).0.this\.\ExponentSizeSize\ := to_unsigned(4, 8);
                        \UnumEnvironment::.ctor(Byte,Byte).0.this\.\FractionSizeSize\ := to_unsigned(8, 8);
                        -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.UnumHelper::SegmentSizeSizeToSegmentSize(System.Byte)
                        \UnumEnvironment::.ctor(Byte,Byte).0.UnumHelper::SegmentSizeSizeToSegmentSize(Byte).segmentSizeSize.parameter.Out.0\ <= to_unsigned(4, 8);
                        \UnumEnvironment::.ctor(Byte,Byte).0.UnumHelper::SegmentSizeSizeToSegmentSize(Byte)._Started.0\ <= true;
                        \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.UnumHelper::SegmentSizeSizeToSegmentSize(System.Byte)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.UnumHelper::SegmentSizeSizeToSegmentSize(Byte)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.UnumHelper::SegmentSizeSizeToSegmentSize(Byte)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.UnumHelper::SegmentSizeSizeToSegmentSize(Byte)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.return.0\ := \UnumEnvironment::.ctor(Byte,Byte).0.UnumHelper::SegmentSizeSizeToSegmentSize(Byte).return.0\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\ExponentSizeMax\ := resize(\UnumEnvironment::.ctor(Byte,Byte).0.return.0\, 8);
                            -- The last invocation for the target state machine just finished, so need to start the next one in a later state.
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_4\ => 
                        -- This state was just added to leave time for the invocation proxy to register that the previous invocation finished.
                        \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_5\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_5\ => 
                        -- Starting state machine invocation for the following method: System.UInt16 Lombiq.Unum.UnumHelper::SegmentSizeSizeToSegmentSize(System.Byte)
                        \UnumEnvironment::.ctor(Byte,Byte).0.UnumHelper::SegmentSizeSizeToSegmentSize(Byte).segmentSizeSize.parameter.Out.0\ <= to_unsigned(8, 8);
                        \UnumEnvironment::.ctor(Byte,Byte).0.UnumHelper::SegmentSizeSizeToSegmentSize(Byte)._Started.0\ <= true;
                        \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_6\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_6\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.UInt16 Lombiq.Unum.UnumHelper::SegmentSizeSizeToSegmentSize(System.Byte)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.UnumHelper::SegmentSizeSizeToSegmentSize(Byte)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.UnumHelper::SegmentSizeSizeToSegmentSize(Byte)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.UnumHelper::SegmentSizeSizeToSegmentSize(Byte)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.return.1\ := \UnumEnvironment::.ctor(Byte,Byte).0.UnumHelper::SegmentSizeSizeToSegmentSize(Byte).return.0\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\FractionSizeMax\ := \UnumEnvironment::.ctor(Byte,Byte).0.return.1\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\UnumTagSize\ := to_unsigned(13, 8);
                            \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.0\ := resize(to_unsigned(1, 8) + \UnumEnvironment::.ctor(Byte,Byte).0.this\.\ExponentSizeMax\, 16);
                            \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.1\ := resize((\UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.0\) + \UnumEnvironment::.ctor(Byte,Byte).0.this\.\FractionSizeMax\, 16);
                            \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.2\ := \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.1\ + to_unsigned(13, 16);
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\Size\ := \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.2\;
                            -- Initializing record fields to their defaults.
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\EmptyBitMask\.\IsNull\ := false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\EmptyBitMask\.\Size\ := to_unsigned(0, 16);
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\EmptyBitMask\.\SegmentCount\ := to_unsigned(0, 16);
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\EmptyBitMask\.\Segments\ := (others => to_unsigned(0, 32));
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\EmptyBitMask\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\Size\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\ <= False;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= true;
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_7\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\EmptyBitMask\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\;
                            -- Initializing record fields to their defaults.
                            \UnumEnvironment::.ctor(Byte,Byte).0.objecta4c70e00f2ec2975ffd03b87442e75fb219dd43f089d457c217e1f67cffbf4a0\.\IsNull\ := false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.objecta4c70e00f2ec2975ffd03b87442e75fb219dd43f089d457c217e1f67cffbf4a0\.\Size\ := to_unsigned(0, 16);
                            \UnumEnvironment::.ctor(Byte,Byte).0.objecta4c70e00f2ec2975ffd03b87442e75fb219dd43f089d457c217e1f67cffbf4a0\.\SegmentCount\ := to_unsigned(0, 16);
                            \UnumEnvironment::.ctor(Byte,Byte).0.objecta4c70e00f2ec2975ffd03b87442e75fb219dd43f089d457c217e1f67cffbf4a0\.\Segments\ := (others => to_unsigned(0, 32));
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.objecta4c70e00f2ec2975ffd03b87442e75fb219dd43f089d457c217e1f67cffbf4a0\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\Size\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\ <= False;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= true;
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_8\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.objecta4c70e00f2ec2975ffd03b87442e75fb219dd43f089d457c217e1f67cffbf4a0\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetOne(System.UInt16)
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).this.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.objecta4c70e00f2ec2975ffd03b87442e75fb219dd43f089d457c217e1f67cffbf4a0\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).index.parameter.Out.0\ <= to_unsigned(12, 16);
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Started.0\ <= true;
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_9\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_9\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetOne(System.UInt16)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.return.2\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).return.0\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\UncertaintyBitMask\ := \UnumEnvironment::.ctor(Byte,Byte).0.return.2\;
                            -- Initializing record fields to their defaults.
                            \UnumEnvironment::.ctor(Byte,Byte).0.object1af8c7e1413e2da44291e3b4786150cb23fed68c0d70afe08a2e21d86ea1dbf3\.\IsNull\ := false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.object1af8c7e1413e2da44291e3b4786150cb23fed68c0d70afe08a2e21d86ea1dbf3\.\Size\ := to_unsigned(0, 16);
                            \UnumEnvironment::.ctor(Byte,Byte).0.object1af8c7e1413e2da44291e3b4786150cb23fed68c0d70afe08a2e21d86ea1dbf3\.\SegmentCount\ := to_unsigned(0, 16);
                            \UnumEnvironment::.ctor(Byte,Byte).0.object1af8c7e1413e2da44291e3b4786150cb23fed68c0d70afe08a2e21d86ea1dbf3\.\Segments\ := (others => to_unsigned(0, 32));
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.object1af8c7e1413e2da44291e3b4786150cb23fed68c0d70afe08a2e21d86ea1dbf3\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\Size\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\ <= False;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= true;
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_10\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_10\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.object1af8c7e1413e2da44291e3b4786150cb23fed68c0d70afe08a2e21d86ea1dbf3\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\;
                            -- The last invocation for the target state machine finished in the previous state, so need to start the next one in the next state.
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_11\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_11\ => 
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetOne(System.UInt16)
                        \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).this.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.object1af8c7e1413e2da44291e3b4786150cb23fed68c0d70afe08a2e21d86ea1dbf3\;
                        \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).index.parameter.Out.0\ <= to_unsigned(8, 16);
                        \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Started.0\ <= true;
                        \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_12\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_12\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetOne(System.UInt16)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.return.3\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,System.UInt32)
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).left.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.return.3\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).right.parameter.Out.0\ <= to_unsigned(1, 32);
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ <= true;
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_13\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_13\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,System.UInt32)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.return.4\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).return.0\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\FractionSizeMask\ := \UnumEnvironment::.ctor(Byte,Byte).0.return.4\;
                            -- The last invocation for the target state machine just finished, so need to start the next one in a later state.
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_14\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_14\ => 
                        -- This state was just added to leave time for the invocation proxy to register that the previous invocation finished.
                        \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_15\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_15\ => 
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,System.UInt32)
                        \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).left.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\UncertaintyBitMask\;
                        \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).right.parameter.Out.0\ <= to_unsigned(1, 32);
                        \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ <= true;
                        \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_16\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_16\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,System.UInt32)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.return.5\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask).left.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.return.5\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask).right.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\FractionSizeMask\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ <= true;
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_17\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_17\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.return.6\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask).return.0\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\ExponentSizeMask\ := \UnumEnvironment::.ctor(Byte,Byte).0.return.6\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseOr(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_BitwiseOr(BitMask,BitMask).left.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\ExponentSizeMask\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_BitwiseOr(BitMask,BitMask).right.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\FractionSizeMask\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_BitwiseOr(BitMask,BitMask)._Started.0\ <= true;
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_18\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_18\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseOr(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_BitwiseOr(BitMask,BitMask)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_BitwiseOr(BitMask,BitMask)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_BitwiseOr(BitMask,BitMask)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.return.7\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_BitwiseOr(BitMask,BitMask).return.0\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\ExponentAndFractionSizeMask\ := \UnumEnvironment::.ctor(Byte,Byte).0.return.7\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask).left.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\UncertaintyBitMask\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask).right.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\ExponentAndFractionSizeMask\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= true;
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_19\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_19\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.return.8\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask).return.0\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\UnumTagMask\ := \UnumEnvironment::.ctor(Byte,Byte).0.return.8\;
                            -- Initializing record fields to their defaults.
                            \UnumEnvironment::.ctor(Byte,Byte).0.object7f34fefc400743c5659b915282ee58959b74703089d82e84e8d6c948e4b443d7\.\IsNull\ := false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.object7f34fefc400743c5659b915282ee58959b74703089d82e84e8d6c948e4b443d7\.\Size\ := to_unsigned(0, 16);
                            \UnumEnvironment::.ctor(Byte,Byte).0.object7f34fefc400743c5659b915282ee58959b74703089d82e84e8d6c948e4b443d7\.\SegmentCount\ := to_unsigned(0, 16);
                            \UnumEnvironment::.ctor(Byte,Byte).0.object7f34fefc400743c5659b915282ee58959b74703089d82e84e8d6c948e4b443d7\.\Segments\ := (others => to_unsigned(0, 32));
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.object7f34fefc400743c5659b915282ee58959b74703089d82e84e8d6c948e4b443d7\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\Size\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\ <= False;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= true;
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_20\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_20\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.object7f34fefc400743c5659b915282ee58959b74703089d82e84e8d6c948e4b443d7\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.3\ := \UnumEnvironment::.ctor(Byte,Byte).0.this\.\Size\ - to_unsigned(1, 16);
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetOne(System.UInt16)
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).this.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.object7f34fefc400743c5659b915282ee58959b74703089d82e84e8d6c948e4b443d7\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).index.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.3\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Started.0\ <= true;
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_21\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_21\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetOne(System.UInt16)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.return.9\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).return.0\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\SignBitMask\ := \UnumEnvironment::.ctor(Byte,Byte).0.return.9\;
                            -- Initializing record fields to their defaults.
                            \UnumEnvironment::.ctor(Byte,Byte).0.objecte438b2d1e01c6422c441d4244fd563f19ddf9cd04a02503bb4f07fbb1fcf4864\.\IsNull\ := false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.objecte438b2d1e01c6422c441d4244fd563f19ddf9cd04a02503bb4f07fbb1fcf4864\.\Size\ := to_unsigned(0, 16);
                            \UnumEnvironment::.ctor(Byte,Byte).0.objecte438b2d1e01c6422c441d4244fd563f19ddf9cd04a02503bb4f07fbb1fcf4864\.\SegmentCount\ := to_unsigned(0, 16);
                            \UnumEnvironment::.ctor(Byte,Byte).0.objecte438b2d1e01c6422c441d4244fd563f19ddf9cd04a02503bb4f07fbb1fcf4864\.\Segments\ := (others => to_unsigned(0, 32));
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.objecte438b2d1e01c6422c441d4244fd563f19ddf9cd04a02503bb4f07fbb1fcf4864\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\Size\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\ <= False;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= true;
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_22\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_22\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.objecte438b2d1e01c6422c441d4244fd563f19ddf9cd04a02503bb4f07fbb1fcf4864\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\;
                            -- The last invocation for the target state machine finished in the previous state, so need to start the next one in the next state.
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_23\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_23\ => 
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetOne(System.UInt16)
                        \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).this.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.objecte438b2d1e01c6422c441d4244fd563f19ddf9cd04a02503bb4f07fbb1fcf4864\;
                        \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).index.parameter.Out.0\ <= to_unsigned(13, 16);
                        \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Started.0\ <= true;
                        \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_24\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_24\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetOne(System.UInt16)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.return.10\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).return.0\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\ULP\ := \UnumEnvironment::.ctor(Byte,Byte).0.return.10\;
                            -- Initializing record fields to their defaults.
                            \UnumEnvironment::.ctor(Byte,Byte).0.object479fe084fa4366b617a7eeccf1cdebf1ed267e764cb62ef8fe9d94f131cbeab7\.\IsNull\ := false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.object479fe084fa4366b617a7eeccf1cdebf1ed267e764cb62ef8fe9d94f131cbeab7\.\Size\ := to_unsigned(0, 16);
                            \UnumEnvironment::.ctor(Byte,Byte).0.object479fe084fa4366b617a7eeccf1cdebf1ed267e764cb62ef8fe9d94f131cbeab7\.\SegmentCount\ := to_unsigned(0, 16);
                            \UnumEnvironment::.ctor(Byte,Byte).0.object479fe084fa4366b617a7eeccf1cdebf1ed267e764cb62ef8fe9d94f131cbeab7\.\Segments\ := (others => to_unsigned(0, 32));
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.object479fe084fa4366b617a7eeccf1cdebf1ed267e764cb62ef8fe9d94f131cbeab7\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\Size\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\ <= False;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= true;
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_25\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_25\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.object479fe084fa4366b617a7eeccf1cdebf1ed267e764cb62ef8fe9d94f131cbeab7\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.4\ := \UnumEnvironment::.ctor(Byte,Byte).0.this\.\Size\ - to_unsigned(1, 16);
                            -- The last invocation for the target state machine finished in the previous state, so need to start the next one in the next state.
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_26\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_26\ => 
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetOne(System.UInt16)
                        \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).this.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.object479fe084fa4366b617a7eeccf1cdebf1ed267e764cb62ef8fe9d94f131cbeab7\;
                        \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).index.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.4\;
                        \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Started.0\ <= true;
                        \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_27\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_27\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetOne(System.UInt16)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.return.11\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,System.UInt32)
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).left.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.return.11\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).right.parameter.Out.0\ <= to_unsigned(1, 32);
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ <= true;
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_28\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_28\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,System.UInt32)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.return.12\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask).left.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.return.12\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask).right.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\UncertaintyBitMask\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ <= true;
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_29\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_29\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.return.13\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask).return.0\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\PositiveInfinity\ := \UnumEnvironment::.ctor(Byte,Byte).0.return.13\;
                            -- Initializing record fields to their defaults.
                            \UnumEnvironment::.ctor(Byte,Byte).0.objectf4f045d4d2f66a18d2b9627940ae5ecef55676a7cd16373be4c2abd2bc60efc2\.\IsNull\ := false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.objectf4f045d4d2f66a18d2b9627940ae5ecef55676a7cd16373be4c2abd2bc60efc2\.\Size\ := to_unsigned(0, 16);
                            \UnumEnvironment::.ctor(Byte,Byte).0.objectf4f045d4d2f66a18d2b9627940ae5ecef55676a7cd16373be4c2abd2bc60efc2\.\SegmentCount\ := to_unsigned(0, 16);
                            \UnumEnvironment::.ctor(Byte,Byte).0.objectf4f045d4d2f66a18d2b9627940ae5ecef55676a7cd16373be4c2abd2bc60efc2\.\Segments\ := (others => to_unsigned(0, 32));
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.objectf4f045d4d2f66a18d2b9627940ae5ecef55676a7cd16373be4c2abd2bc60efc2\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\Size\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\ <= False;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= true;
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_30\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_30\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.objectf4f045d4d2f66a18d2b9627940ae5ecef55676a7cd16373be4c2abd2bc60efc2\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.5\ := \UnumEnvironment::.ctor(Byte,Byte).0.this\.\Size\ - to_unsigned(1, 16);
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetOne(System.UInt16)
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).this.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.objectf4f045d4d2f66a18d2b9627940ae5ecef55676a7cd16373be4c2abd2bc60efc2\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).index.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.5\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Started.0\ <= true;
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_31\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_31\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetOne(System.UInt16)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.return.14\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).return.0\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask).left.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.return.14\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask).right.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\PositiveInfinity\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= true;
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_32\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_32\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.return.15\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask).return.0\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\NegativeInfinity\ := \UnumEnvironment::.ctor(Byte,Byte).0.return.15\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask).left.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\PositiveInfinity\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask).right.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\ULP\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ <= true;
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_33\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_33\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.return.16\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask).return.0\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\LargestPositive\ := \UnumEnvironment::.ctor(Byte,Byte).0.return.16\;
                            -- The last invocation for the target state machine finished in the previous state, so need to start the next one in the next state.
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_34\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_34\ => 
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask).left.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\ExponentAndFractionSizeMask\;
                        \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask).right.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\ULP\;
                        \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= true;
                        \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_35\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_35\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.return.17\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask).return.0\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\SmallestPositive\ := \UnumEnvironment::.ctor(Byte,Byte).0.return.17\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask).left.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\NegativeInfinity\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask).right.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\ULP\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ <= true;
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_36\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_36\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.return.18\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask).return.0\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\LargestNegative\ := \UnumEnvironment::.ctor(Byte,Byte).0.return.18\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.6\ := resize(signed(\UnumEnvironment::.ctor(Byte,Byte).0.this\.\Size\ - to_unsigned(1, 16)), 32);
                            \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.7\ := resize(shift_left(to_unsigned(1, 32), to_integer((\UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.6\))), 32);
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,System.UInt32)
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,UInt32).left.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\LargestPositive\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.binaryOperationResult.7\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ <= true;
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_37\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_37\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,System.UInt32)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.return.19\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,UInt32).return.0\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\MinRealU\ := \UnumEnvironment::.ctor(Byte,Byte).0.return.19\;
                            -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask).left.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\PositiveInfinity\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask).right.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\UncertaintyBitMask\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= true;
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_38\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_38\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.return.20\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask).return.0\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\QuietNotANumber\ := \UnumEnvironment::.ctor(Byte,Byte).0.return.20\;
                            -- The last invocation for the target state machine just finished, so need to start the next one in a later state.
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_39\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_39\ => 
                        -- This state was just added to leave time for the invocation proxy to register that the previous invocation finished.
                        \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_40\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_40\ => 
                        -- Starting state machine invocation for the following method: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask).left.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\NegativeInfinity\;
                        \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask).right.parameter.Out.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this\.\UncertaintyBitMask\;
                        \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= true;
                        \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_41\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnumEnvironment::.ctor(Byte,Byte).0._State_41\ => 
                        -- Waiting for the state machine invocation of the following method to finish: Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask)
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ = \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ <= false;
                            \UnumEnvironment::.ctor(Byte,Byte).0.return.21\ := \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask).return.0\;
                            \UnumEnvironment::.ctor(Byte,Byte).0.this\.\SignalingNotANumber\ := \UnumEnvironment::.ctor(Byte,Byte).0.return.21\;
                            \UnumEnvironment::.ctor(Byte,Byte).0._State\ := \UnumEnvironment::.ctor(Byte,Byte).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Lombiq.Unum.UnumEnvironment::.ctor(System.Byte,System.Byte).0 state machine end


    -- System.Void Hast::ExternalInvocationProxy() start
    \Finished\ <= \FinishedInternal\;
    \Hast::ExternalInvocationProxy()\: process (\Clock\) 
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \FinishedInternal\ <= false;
                \Hast::ExternalInvocationProxy().UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory)._Started.0\ <= false;
            else 
                if (\Started\ = true and \FinishedInternal\ = false) then 
                    -- Starting the state machine corresponding to the given member ID.
                    case \MemberId\ is 
                        when 0 => 
                            if (\Hast::ExternalInvocationProxy().UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory)._Started.0\ = \Hast::ExternalInvocationProxy().UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when others => 
                            null;
                    end case;
                else 
                    -- Waiting for Started to be pulled back to zero that signals the framework noting the finish.
                    if (\Started\ = false and \FinishedInternal\ = true) then 
                        \FinishedInternal\ <= false;
                    end if;
                end if;
            end if;
        end if;
    end process;
    -- System.Void Hast::ExternalInvocationProxy() end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.UnumEnvironment Hast.Samples.SampleAssembly.UnumCalculator::EnvironmentFactory() start
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.UnumCalculator::CalculateSumOfPowersofTwo(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 (#0):
    \UnumCalculator::EnvironmentFactory().0._Started\ <= \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.UnumCalculator::EnvironmentFactory()._Started.0\;
    \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.UnumCalculator::EnvironmentFactory()._Finished.0\ <= \UnumCalculator::EnvironmentFactory().0._Finished\;
    \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.UnumCalculator::EnvironmentFactory().return.0\ <= \UnumCalculator::EnvironmentFactory().0.return\;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.UnumEnvironment Hast.Samples.SampleAssembly.UnumCalculator::EnvironmentFactory() end


    -- System.Void Hast::InternalInvocationProxy().System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.Int32) start
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.UnumCalculator::CalculateSumOfPowersofTwo(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 (#0):
    \Unum::.ctor(UnumEnvironment,Int32).0._Started\ <= \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32)._Started.0\;
    \Unum::.ctor(UnumEnvironment,Int32).0.this.parameter.In\ <= \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32).this.parameter.Out.0\;
    \Unum::.ctor(UnumEnvironment,Int32).0.environment.parameter.In\ <= \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32).environment.parameter.Out.0\;
    \Unum::.ctor(UnumEnvironment,Int32).0.value.parameter.In\ <= \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32).value.parameter.Out.0\;
    \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32)._Finished.0\ <= \Unum::.ctor(UnumEnvironment,Int32).0._Finished\;
    \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32).this.parameter.In.0\ <= \Unum::.ctor(UnumEnvironment,Int32).0.this.parameter.Out\;
    \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::.ctor(UnumEnvironment,Int32).environment.parameter.In.0\ <= \Unum::.ctor(UnumEnvironment,Int32).0.environment.parameter.Out\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.Int32) end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.Unum Lombiq.Unum.Unum::op_Addition(Lombiq.Unum.Unum,Lombiq.Unum.Unum) start
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.UnumCalculator::CalculateSumOfPowersofTwo(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 (#0):
    \Unum::op_Addition(Unum,Unum).0._Started\ <= \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum)._Started.0\;
    \Unum::op_Addition(Unum,Unum).0.left.parameter.In\ <= \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum).left.parameter.Out.0\;
    \Unum::op_Addition(Unum,Unum).0.right.parameter.In\ <= \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum).right.parameter.Out.0\;
    \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum)._Finished.0\ <= \Unum::op_Addition(Unum,Unum).0._Finished\;
    \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::op_Addition(Unum,Unum).return.0\ <= \Unum::op_Addition(Unum,Unum).0.return\;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.Unum Lombiq.Unum.Unum::op_Addition(Lombiq.Unum.Unum,Lombiq.Unum.Unum) end


    -- System.Void Hast::InternalInvocationProxy().System.UInt32[] Lombiq.Unum.Unum::FractionToUintArray() start
    -- Signal connections for System.Void Hast.Samples.SampleAssembly.UnumCalculator::CalculateSumOfPowersofTwo(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory).0 (#0):
    \Unum::FractionToUintArray().0._Started\ <= \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::FractionToUintArray()._Started.0\;
    \Unum::FractionToUintArray().0.this.parameter.In\ <= \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::FractionToUintArray().this.parameter.Out.0\;
    \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::FractionToUintArray()._Finished.0\ <= \Unum::FractionToUintArray().0._Finished\;
    \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.Unum::FractionToUintArray().return.0\ <= \Unum::FractionToUintArray().0.return\;
    -- System.Void Hast::InternalInvocationProxy().System.UInt32[] Lombiq.Unum.Unum::FractionToUintArray() end


    -- System.Void Hast::InternalInvocationProxy().System.Void Lombiq.Unum.UnumEnvironment::.ctor(System.Byte,System.Byte) start
    -- Signal connections for Lombiq.Unum.UnumEnvironment Hast.Samples.SampleAssembly.UnumCalculator::EnvironmentFactory().0 (#0):
    \UnumEnvironment::.ctor(Byte,Byte).0._Started\ <= \UnumCalculator::EnvironmentFactory().0.UnumEnvironment::.ctor(Byte,Byte)._Started.0\;
    \UnumEnvironment::.ctor(Byte,Byte).0.this.parameter.In\ <= \UnumCalculator::EnvironmentFactory().0.UnumEnvironment::.ctor(Byte,Byte).this.parameter.Out.0\;
    \UnumEnvironment::.ctor(Byte,Byte).0.exponentSizeSize.parameter.In\ <= \UnumCalculator::EnvironmentFactory().0.UnumEnvironment::.ctor(Byte,Byte).exponentSizeSize.parameter.Out.0\;
    \UnumEnvironment::.ctor(Byte,Byte).0.fractionSizeSize.parameter.In\ <= \UnumCalculator::EnvironmentFactory().0.UnumEnvironment::.ctor(Byte,Byte).fractionSizeSize.parameter.Out.0\;
    \UnumCalculator::EnvironmentFactory().0.UnumEnvironment::.ctor(Byte,Byte)._Finished.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0._Finished\;
    \UnumCalculator::EnvironmentFactory().0.UnumEnvironment::.ctor(Byte,Byte).this.parameter.In.0\ <= \UnumEnvironment::.ctor(Byte,Byte).0.this.parameter.Out\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Lombiq.Unum.UnumEnvironment::.ctor(System.Byte,System.Byte) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16) start
    \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::FromImmutableArray(UInt32[],UInt16).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::FromImmutableArray(UInt32[],UInt16).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Addition(BitMask,UInt32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Addition(BitMask,UInt32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Subtraction(BitMask,UInt32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Subtraction(BitMask,UInt32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Addition(BitMask,BitMask).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Addition(BitMask,BitMask).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Subtraction(BitMask,BitMask).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Subtraction(BitMask,BitMask).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_BitwiseOr(BitMask,BitMask).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_BitwiseOr(BitMask,BitMask).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_BitwiseAnd(BitMask,BitMask).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_BitwiseAnd(BitMask,BitMask).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_RightShift(BitMask,Int32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_RightShift(BitMask,Int32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_LeftShift(BitMask,Int32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_LeftShift(BitMask,Int32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::FractionMask().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::FractionMask().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::ExponentMask().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::ExponentMask().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::FromImmutableArray(UInt32[],UInt16).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::FromImmutableArray(UInt32[],UInt16).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Addition(BitMask,UInt32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Addition(BitMask,UInt32).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Subtraction(BitMask,UInt32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Subtraction(BitMask,UInt32).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Addition(BitMask,BitMask).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Addition(BitMask,BitMask).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Subtraction(BitMask,BitMask).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Subtraction(BitMask,BitMask).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_BitwiseOr(BitMask,BitMask).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_BitwiseOr(BitMask,BitMask).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_BitwiseAnd(BitMask,BitMask).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_BitwiseAnd(BitMask,BitMask).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_RightShift(BitMask,Int32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_RightShift(BitMask,Int32).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_LeftShift(BitMask,Int32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_LeftShift(BitMask,Int32).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::FractionMask().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::FractionMask().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::ExponentMask().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::ExponentMask().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningState.0\ := WaitingForStarted;
                \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.BitMask::FromImmutableArray(System.UInt32[],System.UInt16).0
                case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::FromImmutableArray(UInt32[],UInt16).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\) then 
                            \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::FromImmutableArray(UInt32[],UInt16).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::FromImmutableArray(UInt32[],UInt16).0.runningIndex.0\ := 0;
                            \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= true;
                            \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.In\ <= \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.In\ <= \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.size.parameter.In\ <= \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::FromImmutableArray(UInt32[],UInt16).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::.ctor(UInt32[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::FromImmutableArray(UInt32[],UInt16).0.runningState.0\ := AfterFinished;
                                    \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= true;
                                    \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= false;
                                    \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.Out\;
                                    \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::FromImmutableArray(UInt32[],UInt16).0.runningState.0\ := WaitingForStarted;
                            \BitMask::FromImmutableArray(UInt32[],UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,System.UInt32).0
                case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Addition(BitMask,UInt32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\) then 
                            \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Addition(BitMask,UInt32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Addition(BitMask,UInt32).0.runningIndex.0\ := 0;
                            \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= true;
                            \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.In\ <= \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.In\ <= \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.size.parameter.In\ <= \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Addition(BitMask,UInt32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::.ctor(UInt32[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Addition(BitMask,UInt32).0.runningState.0\ := AfterFinished;
                                    \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= true;
                                    \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= false;
                                    \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.Out\;
                                    \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Addition(BitMask,UInt32).0.runningState.0\ := WaitingForStarted;
                            \BitMask::op_Addition(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,System.UInt32).0
                case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Subtraction(BitMask,UInt32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\) then 
                            \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Subtraction(BitMask,UInt32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Subtraction(BitMask,UInt32).0.runningIndex.0\ := 0;
                            \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= true;
                            \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.In\ <= \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.In\ <= \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.size.parameter.In\ <= \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Subtraction(BitMask,UInt32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::.ctor(UInt32[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Subtraction(BitMask,UInt32).0.runningState.0\ := AfterFinished;
                                    \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= true;
                                    \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= false;
                                    \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.Out\;
                                    \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Subtraction(BitMask,UInt32).0.runningState.0\ := WaitingForStarted;
                            \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0
                case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Addition(BitMask,BitMask).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\) then 
                            \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Addition(BitMask,BitMask).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Addition(BitMask,BitMask).0.runningIndex.0\ := 0;
                            \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= true;
                            \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.In\ <= \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.In\ <= \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.size.parameter.In\ <= \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Addition(BitMask,BitMask).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::.ctor(UInt32[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Addition(BitMask,BitMask).0.runningState.0\ := AfterFinished;
                                    \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= true;
                                    \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= false;
                                    \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.Out\;
                                    \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Addition(BitMask,BitMask).0.runningState.0\ := WaitingForStarted;
                            \BitMask::op_Addition(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0
                case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Subtraction(BitMask,BitMask).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\) then 
                            \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Subtraction(BitMask,BitMask).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Subtraction(BitMask,BitMask).0.runningIndex.0\ := 0;
                            \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= true;
                            \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.In\ <= \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.In\ <= \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.size.parameter.In\ <= \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Subtraction(BitMask,BitMask).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::.ctor(UInt32[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Subtraction(BitMask,BitMask).0.runningState.0\ := AfterFinished;
                                    \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= true;
                                    \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= false;
                                    \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.Out\;
                                    \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_Subtraction(BitMask,BitMask).0.runningState.0\ := WaitingForStarted;
                            \BitMask::op_Subtraction(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseOr(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0
                case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_BitwiseOr(BitMask,BitMask).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\) then 
                            \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_BitwiseOr(BitMask,BitMask).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_BitwiseOr(BitMask,BitMask).0.runningIndex.0\ := 0;
                            \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= true;
                            \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.In\ <= \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.In\ <= \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.size.parameter.In\ <= \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_BitwiseOr(BitMask,BitMask).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::.ctor(UInt32[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_BitwiseOr(BitMask,BitMask).0.runningState.0\ := AfterFinished;
                                    \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= true;
                                    \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= false;
                                    \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.Out\;
                                    \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_BitwiseOr(BitMask,BitMask).0.runningState.0\ := WaitingForStarted;
                            \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseAnd(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0
                case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_BitwiseAnd(BitMask,BitMask).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\) then 
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_BitwiseAnd(BitMask,BitMask).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_BitwiseAnd(BitMask,BitMask).0.runningIndex.0\ := 0;
                            \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= true;
                            \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.In\ <= \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.In\ <= \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.size.parameter.In\ <= \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_BitwiseAnd(BitMask,BitMask).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::.ctor(UInt32[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_BitwiseAnd(BitMask,BitMask).0.runningState.0\ := AfterFinished;
                                    \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= true;
                                    \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= false;
                                    \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.Out\;
                                    \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_BitwiseAnd(BitMask,BitMask).0.runningState.0\ := WaitingForStarted;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_RightShift(Lombiq.Unum.BitMask,System.Int32).0
                case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_RightShift(BitMask,Int32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\) then 
                            \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_RightShift(BitMask,Int32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_RightShift(BitMask,Int32).0.runningIndex.0\ := 0;
                            \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= true;
                            \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.In\ <= \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.In\ <= \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.size.parameter.In\ <= \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_RightShift(BitMask,Int32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::.ctor(UInt32[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_RightShift(BitMask,Int32).0.runningState.0\ := AfterFinished;
                                    \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= true;
                                    \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= false;
                                    \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.Out\;
                                    \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_RightShift(BitMask,Int32).0.runningState.0\ := WaitingForStarted;
                            \BitMask::op_RightShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32).0
                case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_LeftShift(BitMask,Int32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\) then 
                            \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_LeftShift(BitMask,Int32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_LeftShift(BitMask,Int32).0.runningIndex.0\ := 0;
                            \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= true;
                            \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.In\ <= \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.In\ <= \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.size.parameter.In\ <= \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_LeftShift(BitMask,Int32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::.ctor(UInt32[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_LeftShift(BitMask,Int32).0.runningState.0\ := AfterFinished;
                                    \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= true;
                                    \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= false;
                                    \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.Out\;
                                    \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).BitMask::op_LeftShift(BitMask,Int32).0.runningState.0\ := WaitingForStarted;
                            \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.UInt32[],System.Boolean).0
                case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ := 0;
                            \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= true;
                            \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.In\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.In\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.size.parameter.In\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::.ctor(UInt32[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := AfterFinished;
                                    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= true;
                                    \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= false;
                                    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.Out\;
                                    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForStarted;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::SetUnumBits(System.Boolean,Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean,System.Byte,System.UInt16).0
                case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\) then 
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\ := 0;
                            \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= true;
                            \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.In\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.In\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.size.parameter.In\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::.ctor(UInt32[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := AfterFinished;
                                    \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= true;
                                    \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= false;
                                    \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.Out\;
                                    \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := WaitingForStarted;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionMask().0
                case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::FractionMask().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16)._Started.0\) then 
                            \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::FractionMask().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::FractionMask().0.runningIndex.0\ := 0;
                            \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= true;
                            \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.In\ <= \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.In\ <= \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.size.parameter.In\ <= \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::FractionMask().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::.ctor(UInt32[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::FractionMask().0.runningState.0\ := AfterFinished;
                                    \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= true;
                                    \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= false;
                                    \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.Out\;
                                    \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::FractionMask().0.runningState.0\ := WaitingForStarted;
                            \Unum::FractionMask().0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentMask().0
                case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::ExponentMask().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16)._Started.0\) then 
                            \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::ExponentMask().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::ExponentMask().0.runningIndex.0\ := 0;
                            \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= true;
                            \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.In\ <= \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.In\ <= \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.size.parameter.In\ <= \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::ExponentMask().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::.ctor(UInt32[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::ExponentMask().0.runningState.0\ := AfterFinished;
                                    \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= true;
                                    \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= false;
                                    \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.Out\;
                                    \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::ExponentMask().0.runningState.0\ := WaitingForStarted;
                            \Unum::ExponentMask().0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentValueToExponentBits(System.Int32,System.Byte).0
                case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\) then 
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningIndex.0\ := 0;
                            \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= true;
                            \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.In\ <= \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.In\ <= \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.Out.0\;
                            \BitMask::.ctor(UInt32[],UInt16).0.size.parameter.In\ <= \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::.ctor(UInt32[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningState.0\ := AfterFinished;
                                    \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= true;
                                    \BitMask::.ctor(UInt32[],UInt16).0._Started\ <= false;
                                    \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16).this.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.this.parameter.Out\;
                                    \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16).segments.parameter.In.0\ <= \BitMask::.ctor(UInt32[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt32[],UInt16).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningState.0\ := WaitingForStarted;
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::.ctor(UInt32[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.Void Lombiq.Unum.BitMask::.ctor(System.UInt32[],System.UInt16) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Lombiq.Unum.BitMask::.ctor(Lombiq.Unum.BitMask) start
    \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::SetOne(UInt16).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::SetOne(UInt16).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::SetZero(UInt16).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::SetZero(UInt16).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::ShiftOutLeastSignificantZeros().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::ShiftOutLeastSignificantZeros().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::SetOne(UInt16).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::SetOne(UInt16).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::SetZero(UInt16).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::SetZero(UInt16).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::ShiftOutLeastSignificantZeros().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::ShiftOutLeastSignificantZeros().0.runningState.0\ := WaitingForStarted;
                \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask)._Finished.0\ <= false;
                \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask)._Finished.0\ <= false;
                \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask)._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetOne(System.UInt16).0
                case \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::SetOne(UInt16).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask)._Started.0\) then 
                            \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::SetOne(UInt16).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::SetOne(UInt16).0.runningIndex.0\ := 0;
                            \BitMask::.ctor(BitMask).0._Started\ <= true;
                            \BitMask::.ctor(BitMask).0.this.parameter.In\ <= \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask).this.parameter.Out.0\;
                            \BitMask::.ctor(BitMask).0.source.parameter.In\ <= \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask).source.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::SetOne(UInt16).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::.ctor(BitMask).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::SetOne(UInt16).0.runningState.0\ := AfterFinished;
                                    \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask)._Finished.0\ <= true;
                                    \BitMask::.ctor(BitMask).0._Started\ <= false;
                                    \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask).this.parameter.In.0\ <= \BitMask::.ctor(BitMask).0.this.parameter.Out\;
                                    \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask).source.parameter.In.0\ <= \BitMask::.ctor(BitMask).0.source.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::SetOne(UInt16).0.runningState.0\ := WaitingForStarted;
                            \BitMask::SetOne(UInt16).0.BitMask::.ctor(BitMask)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetZero(System.UInt16).0
                case \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::SetZero(UInt16).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask)._Started.0\) then 
                            \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::SetZero(UInt16).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::SetZero(UInt16).0.runningIndex.0\ := 0;
                            \BitMask::.ctor(BitMask).0._Started\ <= true;
                            \BitMask::.ctor(BitMask).0.this.parameter.In\ <= \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask).this.parameter.Out.0\;
                            \BitMask::.ctor(BitMask).0.source.parameter.In\ <= \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask).source.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::SetZero(UInt16).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::.ctor(BitMask).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::SetZero(UInt16).0.runningState.0\ := AfterFinished;
                                    \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask)._Finished.0\ <= true;
                                    \BitMask::.ctor(BitMask).0._Started\ <= false;
                                    \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask).this.parameter.In.0\ <= \BitMask::.ctor(BitMask).0.this.parameter.Out\;
                                    \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask).source.parameter.In.0\ <= \BitMask::.ctor(BitMask).0.source.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::SetZero(UInt16).0.runningState.0\ := WaitingForStarted;
                            \BitMask::SetZero(UInt16).0.BitMask::.ctor(BitMask)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.BitMask::ShiftOutLeastSignificantZeros().0
                case \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::ShiftOutLeastSignificantZeros().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask)._Started.0\) then 
                            \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::ShiftOutLeastSignificantZeros().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::ShiftOutLeastSignificantZeros().0.runningIndex.0\ := 0;
                            \BitMask::.ctor(BitMask).0._Started\ <= true;
                            \BitMask::.ctor(BitMask).0.this.parameter.In\ <= \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask).this.parameter.Out.0\;
                            \BitMask::.ctor(BitMask).0.source.parameter.In\ <= \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask).source.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::ShiftOutLeastSignificantZeros().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::.ctor(BitMask).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::ShiftOutLeastSignificantZeros().0.runningState.0\ := AfterFinished;
                                    \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask)._Finished.0\ <= true;
                                    \BitMask::.ctor(BitMask).0._Started\ <= false;
                                    \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask).this.parameter.In.0\ <= \BitMask::.ctor(BitMask).0.this.parameter.Out\;
                                    \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask).source.parameter.In.0\ <= \BitMask::.ctor(BitMask).0.source.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::.ctor(BitMask).BitMask::ShiftOutLeastSignificantZeros().0.runningState.0\ := WaitingForStarted;
                            \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::.ctor(BitMask)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.Void Lombiq.Unum.BitMask::.ctor(Lombiq.Unum.BitMask) end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::FromImmutableArray(System.UInt32[],System.UInt16) start
    \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).BitMask::SetOne(UInt16).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).BitMask::SetOne(UInt16).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).BitMask::SetZero(UInt16).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).BitMask::SetZero(UInt16).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).Unum::.ctor(UnumEnvironment,BitMask).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).Unum::.ctor(UnumEnvironment,BitMask).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).BitMask::SetOne(UInt16).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).BitMask::SetOne(UInt16).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).BitMask::SetZero(UInt16).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).BitMask::SetZero(UInt16).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).Unum::.ctor(UnumEnvironment,BitMask).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).Unum::.ctor(UnumEnvironment,BitMask).0.runningState.0\ := WaitingForStarted;
                \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Finished.0\ <= false;
                \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Finished.0\ <= false;
                \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetOne(System.UInt16).0
                case \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).BitMask::SetOne(UInt16).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Started.0\) then 
                            \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).BitMask::SetOne(UInt16).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).BitMask::SetOne(UInt16).0.runningIndex.0\ := 0;
                            \BitMask::FromImmutableArray(UInt32[],UInt16).0._Started\ <= true;
                            \BitMask::FromImmutableArray(UInt32[],UInt16).0.segments.parameter.In\ <= \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).segments.parameter.Out.0\;
                            \BitMask::FromImmutableArray(UInt32[],UInt16).0.size.parameter.In\ <= \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).BitMask::SetOne(UInt16).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::FromImmutableArray(UInt32[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).BitMask::SetOne(UInt16).0.runningState.0\ := AfterFinished;
                                    \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Finished.0\ <= true;
                                    \BitMask::FromImmutableArray(UInt32[],UInt16).0._Started\ <= false;
                                    \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).return.0\ <= \BitMask::FromImmutableArray(UInt32[],UInt16).0.return\;
                                    \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).segments.parameter.In.0\ <= \BitMask::FromImmutableArray(UInt32[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).BitMask::SetOne(UInt16).0.runningState.0\ := WaitingForStarted;
                            \BitMask::SetOne(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetZero(System.UInt16).0
                case \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).BitMask::SetZero(UInt16).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Started.0\) then 
                            \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).BitMask::SetZero(UInt16).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).BitMask::SetZero(UInt16).0.runningIndex.0\ := 0;
                            \BitMask::FromImmutableArray(UInt32[],UInt16).0._Started\ <= true;
                            \BitMask::FromImmutableArray(UInt32[],UInt16).0.segments.parameter.In\ <= \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).segments.parameter.Out.0\;
                            \BitMask::FromImmutableArray(UInt32[],UInt16).0.size.parameter.In\ <= \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).BitMask::SetZero(UInt16).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::FromImmutableArray(UInt32[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).BitMask::SetZero(UInt16).0.runningState.0\ := AfterFinished;
                                    \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Finished.0\ <= true;
                                    \BitMask::FromImmutableArray(UInt32[],UInt16).0._Started\ <= false;
                                    \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).return.0\ <= \BitMask::FromImmutableArray(UInt32[],UInt16).0.return\;
                                    \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16).segments.parameter.In.0\ <= \BitMask::FromImmutableArray(UInt32[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).BitMask::SetZero(UInt16).0.runningState.0\ := WaitingForStarted;
                            \BitMask::SetZero(UInt16).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,Lombiq.Unum.BitMask).0
                case \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).Unum::.ctor(UnumEnvironment,BitMask).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Started.0\) then 
                            \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).Unum::.ctor(UnumEnvironment,BitMask).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).Unum::.ctor(UnumEnvironment,BitMask).0.runningIndex.0\ := 0;
                            \BitMask::FromImmutableArray(UInt32[],UInt16).0._Started\ <= true;
                            \BitMask::FromImmutableArray(UInt32[],UInt16).0.segments.parameter.In\ <= \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16).segments.parameter.Out.0\;
                            \BitMask::FromImmutableArray(UInt32[],UInt16).0.size.parameter.In\ <= \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).Unum::.ctor(UnumEnvironment,BitMask).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::FromImmutableArray(UInt32[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).Unum::.ctor(UnumEnvironment,BitMask).0.runningState.0\ := AfterFinished;
                                    \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Finished.0\ <= true;
                                    \BitMask::FromImmutableArray(UInt32[],UInt16).0._Started\ <= false;
                                    \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16).return.0\ <= \BitMask::FromImmutableArray(UInt32[],UInt16).0.return\;
                                    \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16).segments.parameter.In.0\ <= \BitMask::FromImmutableArray(UInt32[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::FromImmutableArray(UInt32[],UInt16).Unum::.ctor(UnumEnvironment,BitMask).0.runningState.0\ := WaitingForStarted;
                            \Unum::.ctor(UnumEnvironment,BitMask).0.BitMask::FromImmutableArray(UInt32[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::FromImmutableArray(System.UInt32[],System.UInt16) end


    -- System.Void Hast::InternalInvocationProxy().System.UInt16 Lombiq.Unum.BitMask::GetLeastSignificantOnePosition() start
    -- Signal connections for Lombiq.Unum.BitMask Lombiq.Unum.BitMask::ShiftOutLeastSignificantZeros().0 (#0):
    \BitMask::GetLeastSignificantOnePosition().0._Started\ <= \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::GetLeastSignificantOnePosition()._Started.0\;
    \BitMask::GetLeastSignificantOnePosition().0.this.parameter.In\ <= \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::GetLeastSignificantOnePosition().this.parameter.Out.0\;
    \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::GetLeastSignificantOnePosition()._Finished.0\ <= \BitMask::GetLeastSignificantOnePosition().0._Finished\;
    \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::GetLeastSignificantOnePosition().return.0\ <= \BitMask::GetLeastSignificantOnePosition().0.return\;
    -- System.Void Hast::InternalInvocationProxy().System.UInt16 Lombiq.Unum.BitMask::GetLeastSignificantOnePosition() end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_RightShift(Lombiq.Unum.BitMask,System.Int32) start
    \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).BitMask::ShiftOutLeastSignificantZeros().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).BitMask::ShiftOutLeastSignificantZeros().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).BitMask::op_LeftShift(BitMask,Int32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).BitMask::op_LeftShift(BitMask,Int32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::ExponentSize().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::ExponentSize().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::Exponent().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::Exponent().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::Fraction().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::Fraction().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).BitMask::ShiftOutLeastSignificantZeros().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).BitMask::ShiftOutLeastSignificantZeros().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).BitMask::op_LeftShift(BitMask,Int32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).BitMask::op_LeftShift(BitMask,Int32).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::ExponentSize().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::ExponentSize().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::Exponent().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::Exponent().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::Fraction().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::Fraction().0.runningState.0\ := WaitingForStarted;
                \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\ <= false;
                \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\ <= false;
                \Unum::ExponentSize().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\ <= false;
                \Unum::Exponent().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\ <= false;
                \Unum::Fraction().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.BitMask::ShiftOutLeastSignificantZeros().0
                case \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).BitMask::ShiftOutLeastSignificantZeros().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\BitMask::ShiftOutLeastSignificantZeros().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\) then 
                            \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).BitMask::ShiftOutLeastSignificantZeros().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).BitMask::ShiftOutLeastSignificantZeros().0.runningIndex.0\ := 0;
                            \BitMask::op_RightShift(BitMask,Int32).0._Started\ <= true;
                            \BitMask::op_RightShift(BitMask,Int32).0.left.parameter.In\ <= \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::op_RightShift(BitMask,Int32).left.parameter.Out.0\;
                            \BitMask::op_RightShift(BitMask,Int32).0.right.parameter.In\ <= \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::op_RightShift(BitMask,Int32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).BitMask::ShiftOutLeastSignificantZeros().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_RightShift(BitMask,Int32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).BitMask::ShiftOutLeastSignificantZeros().0.runningState.0\ := AfterFinished;
                                    \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\ <= true;
                                    \BitMask::op_RightShift(BitMask,Int32).0._Started\ <= false;
                                    \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::op_RightShift(BitMask,Int32).return.0\ <= \BitMask::op_RightShift(BitMask,Int32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\BitMask::ShiftOutLeastSignificantZeros().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).BitMask::ShiftOutLeastSignificantZeros().0.runningState.0\ := WaitingForStarted;
                            \BitMask::ShiftOutLeastSignificantZeros().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32).0
                case \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).BitMask::op_LeftShift(BitMask,Int32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\BitMask::op_LeftShift(BitMask,Int32).0.BitMask::op_RightShift(BitMask,Int32)._Started.0\) then 
                            \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).BitMask::op_LeftShift(BitMask,Int32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).BitMask::op_LeftShift(BitMask,Int32).0.runningIndex.0\ := 0;
                            \BitMask::op_RightShift(BitMask,Int32).0._Started\ <= true;
                            \BitMask::op_RightShift(BitMask,Int32).0.left.parameter.In\ <= \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::op_RightShift(BitMask,Int32).left.parameter.Out.0\;
                            \BitMask::op_RightShift(BitMask,Int32).0.right.parameter.In\ <= \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::op_RightShift(BitMask,Int32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).BitMask::op_LeftShift(BitMask,Int32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_RightShift(BitMask,Int32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).BitMask::op_LeftShift(BitMask,Int32).0.runningState.0\ := AfterFinished;
                                    \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\ <= true;
                                    \BitMask::op_RightShift(BitMask,Int32).0._Started\ <= false;
                                    \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::op_RightShift(BitMask,Int32).return.0\ <= \BitMask::op_RightShift(BitMask,Int32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\BitMask::op_LeftShift(BitMask,Int32).0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).BitMask::op_LeftShift(BitMask,Int32).0.runningState.0\ := WaitingForStarted;
                            \BitMask::op_LeftShift(BitMask,Int32).0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Byte Lombiq.Unum.Unum::ExponentSize().0
                case \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::ExponentSize().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::ExponentSize().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\) then 
                            \Unum::ExponentSize().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::ExponentSize().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::ExponentSize().0.runningIndex.0\ := 0;
                            \BitMask::op_RightShift(BitMask,Int32).0._Started\ <= true;
                            \BitMask::op_RightShift(BitMask,Int32).0.left.parameter.In\ <= \Unum::ExponentSize().0.BitMask::op_RightShift(BitMask,Int32).left.parameter.Out.0\;
                            \BitMask::op_RightShift(BitMask,Int32).0.right.parameter.In\ <= \Unum::ExponentSize().0.BitMask::op_RightShift(BitMask,Int32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::ExponentSize().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_RightShift(BitMask,Int32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::ExponentSize().0.runningState.0\ := AfterFinished;
                                    \Unum::ExponentSize().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\ <= true;
                                    \BitMask::op_RightShift(BitMask,Int32).0._Started\ <= false;
                                    \Unum::ExponentSize().0.BitMask::op_RightShift(BitMask,Int32).return.0\ <= \BitMask::op_RightShift(BitMask,Int32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::ExponentSize().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::ExponentSize().0.runningState.0\ := WaitingForStarted;
                            \Unum::ExponentSize().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::Exponent().0
                case \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::Exponent().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::Exponent().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\) then 
                            \Unum::Exponent().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::Exponent().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::Exponent().0.runningIndex.0\ := 0;
                            \BitMask::op_RightShift(BitMask,Int32).0._Started\ <= true;
                            \BitMask::op_RightShift(BitMask,Int32).0.left.parameter.In\ <= \Unum::Exponent().0.BitMask::op_RightShift(BitMask,Int32).left.parameter.Out.0\;
                            \BitMask::op_RightShift(BitMask,Int32).0.right.parameter.In\ <= \Unum::Exponent().0.BitMask::op_RightShift(BitMask,Int32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::Exponent().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_RightShift(BitMask,Int32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::Exponent().0.runningState.0\ := AfterFinished;
                                    \Unum::Exponent().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\ <= true;
                                    \BitMask::op_RightShift(BitMask,Int32).0._Started\ <= false;
                                    \Unum::Exponent().0.BitMask::op_RightShift(BitMask,Int32).return.0\ <= \BitMask::op_RightShift(BitMask,Int32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::Exponent().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::Exponent().0.runningState.0\ := WaitingForStarted;
                            \Unum::Exponent().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::Fraction().0
                case \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::Fraction().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::Fraction().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\) then 
                            \Unum::Fraction().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::Fraction().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::Fraction().0.runningIndex.0\ := 0;
                            \BitMask::op_RightShift(BitMask,Int32).0._Started\ <= true;
                            \BitMask::op_RightShift(BitMask,Int32).0.left.parameter.In\ <= \Unum::Fraction().0.BitMask::op_RightShift(BitMask,Int32).left.parameter.Out.0\;
                            \BitMask::op_RightShift(BitMask,Int32).0.right.parameter.In\ <= \Unum::Fraction().0.BitMask::op_RightShift(BitMask,Int32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::Fraction().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_RightShift(BitMask,Int32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::Fraction().0.runningState.0\ := AfterFinished;
                                    \Unum::Fraction().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\ <= true;
                                    \BitMask::op_RightShift(BitMask,Int32).0._Started\ <= false;
                                    \Unum::Fraction().0.BitMask::op_RightShift(BitMask,Int32).return.0\ <= \BitMask::op_RightShift(BitMask,Int32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::Fraction().0.BitMask::op_RightShift(BitMask,Int32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_RightShift(BitMask,Int32).Unum::Fraction().0.runningState.0\ := WaitingForStarted;
                            \Unum::Fraction().0.BitMask::op_RightShift(BitMask,Int32)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_RightShift(Lombiq.Unum.BitMask,System.Int32) end


    -- System.Void Hast::InternalInvocationProxy().System.Boolean Lombiq.Unum.BitMask::op_LessThan(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask) start
    -- Signal connections for System.Boolean Lombiq.Unum.BitMask::op_GreaterThanOrEqual(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0 (#0):
    \BitMask::op_LessThan(BitMask,BitMask).0._Started\ <= \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.BitMask::op_LessThan(BitMask,BitMask)._Started.0\;
    \BitMask::op_LessThan(BitMask,BitMask).0.left.parameter.In\ <= \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.BitMask::op_LessThan(BitMask,BitMask).left.parameter.Out.0\;
    \BitMask::op_LessThan(BitMask,BitMask).0.right.parameter.In\ <= \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.BitMask::op_LessThan(BitMask,BitMask).right.parameter.Out.0\;
    \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.BitMask::op_LessThan(BitMask,BitMask)._Finished.0\ <= \BitMask::op_LessThan(BitMask,BitMask).0._Finished\;
    \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.BitMask::op_LessThan(BitMask,BitMask).return.0\ <= \BitMask::op_LessThan(BitMask,BitMask).0.return\;
    -- System.Void Hast::InternalInvocationProxy().System.Boolean Lombiq.Unum.BitMask::op_LessThan(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask) end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask) start
    \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).BitMask::op_Addition(BitMask,UInt32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).BitMask::op_Addition(BitMask,UInt32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::AddExactUnums(Unum,Unum).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).BitMask::op_Addition(BitMask,UInt32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).BitMask::op_Addition(BitMask,UInt32).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := WaitingForStarted;
                \BitMask::op_Addition(BitMask,UInt32).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\ <= false;
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\ <= false;
                \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\ <= false;
                \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,System.UInt32).0
                case \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).BitMask::op_Addition(BitMask,UInt32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\BitMask::op_Addition(BitMask,UInt32).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\) then 
                            \BitMask::op_Addition(BitMask,UInt32).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).BitMask::op_Addition(BitMask,UInt32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).BitMask::op_Addition(BitMask,UInt32).0.runningIndex.0\ := 0;
                            \BitMask::op_Addition(BitMask,BitMask).0._Started\ <= true;
                            \BitMask::op_Addition(BitMask,BitMask).0.left.parameter.In\ <= \BitMask::op_Addition(BitMask,UInt32).0.BitMask::op_Addition(BitMask,BitMask).left.parameter.Out.0\;
                            \BitMask::op_Addition(BitMask,BitMask).0.right.parameter.In\ <= \BitMask::op_Addition(BitMask,UInt32).0.BitMask::op_Addition(BitMask,BitMask).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).BitMask::op_Addition(BitMask,UInt32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Addition(BitMask,BitMask).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).BitMask::op_Addition(BitMask,UInt32).0.runningState.0\ := AfterFinished;
                                    \BitMask::op_Addition(BitMask,UInt32).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\ <= true;
                                    \BitMask::op_Addition(BitMask,BitMask).0._Started\ <= false;
                                    \BitMask::op_Addition(BitMask,UInt32).0.BitMask::op_Addition(BitMask,BitMask).return.0\ <= \BitMask::op_Addition(BitMask,BitMask).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\BitMask::op_Addition(BitMask,UInt32).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).BitMask::op_Addition(BitMask,UInt32).0.runningState.0\ := WaitingForStarted;
                            \BitMask::op_Addition(BitMask,UInt32).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::SetUnumBits(System.Boolean,Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean,System.Byte,System.UInt16).0
                case \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\) then 
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\ := 0;
                            \BitMask::op_Addition(BitMask,BitMask).0._Started\ <= true;
                            \BitMask::op_Addition(BitMask,BitMask).0.left.parameter.In\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask).left.parameter.Out.0\;
                            \BitMask::op_Addition(BitMask,BitMask).0.right.parameter.In\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Addition(BitMask,BitMask).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := AfterFinished;
                                    \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\ <= true;
                                    \BitMask::op_Addition(BitMask,BitMask).0._Started\ <= false;
                                    \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask).return.0\ <= \BitMask::op_Addition(BitMask,BitMask).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := WaitingForStarted;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0
                case \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                            \BitMask::op_Addition(BitMask,BitMask).0._Started\ <= true;
                            \BitMask::op_Addition(BitMask,BitMask).0.left.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_Addition(BitMask,BitMask).left.parameter.Out.0\;
                            \BitMask::op_Addition(BitMask,BitMask).0.right.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_Addition(BitMask,BitMask).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Addition(BitMask,BitMask).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := AfterFinished;
                                    \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\ <= true;
                                    \BitMask::op_Addition(BitMask,BitMask).0._Started\ <= false;
                                    \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_Addition(BitMask,BitMask).return.0\ <= \BitMask::op_Addition(BitMask,BitMask).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::AddAlignedFractions(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean).0
                case \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\) then 
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningIndex.0\ := 0;
                            \BitMask::op_Addition(BitMask,BitMask).0._Started\ <= true;
                            \BitMask::op_Addition(BitMask,BitMask).0.left.parameter.In\ <= \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Addition(BitMask,BitMask).left.parameter.Out.0\;
                            \BitMask::op_Addition(BitMask,BitMask).0.right.parameter.In\ <= \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Addition(BitMask,BitMask).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Addition(BitMask,BitMask).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningState.0\ := AfterFinished;
                                    \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\ <= true;
                                    \BitMask::op_Addition(BitMask,BitMask).0._Started\ <= false;
                                    \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Addition(BitMask,BitMask).return.0\ <= \BitMask::op_Addition(BitMask,BitMask).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningState.0\ := WaitingForStarted;
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Void Lombiq.Unum.UnumEnvironment::.ctor(System.Byte,System.Byte).0
                case \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\ := 0;
                            \BitMask::op_Addition(BitMask,BitMask).0._Started\ <= true;
                            \BitMask::op_Addition(BitMask,BitMask).0.left.parameter.In\ <= \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask).left.parameter.Out.0\;
                            \BitMask::op_Addition(BitMask,BitMask).0.right.parameter.In\ <= \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Addition(BitMask,BitMask).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := AfterFinished;
                                    \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\ <= true;
                                    \BitMask::op_Addition(BitMask,BitMask).0._Started\ <= false;
                                    \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask).return.0\ <= \BitMask::op_Addition(BitMask,BitMask).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,BitMask).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := WaitingForStarted;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,BitMask)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask) end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask) start
    \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).BitMask::op_Subtraction(BitMask,UInt32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).BitMask::op_Subtraction(BitMask,UInt32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).BitMask::op_Subtraction(BitMask,UInt32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).BitMask::op_Subtraction(BitMask,UInt32).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := WaitingForStarted;
                \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::op_Subtraction(BitMask,BitMask)._Finished.0\ <= false;
                \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask)._Finished.0\ <= false;
                \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,System.UInt32).0
                case \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).BitMask::op_Subtraction(BitMask,UInt32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\) then 
                            \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::op_Subtraction(BitMask,BitMask)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).BitMask::op_Subtraction(BitMask,UInt32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).BitMask::op_Subtraction(BitMask,UInt32).0.runningIndex.0\ := 0;
                            \BitMask::op_Subtraction(BitMask,BitMask).0._Started\ <= true;
                            \BitMask::op_Subtraction(BitMask,BitMask).0.left.parameter.In\ <= \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::op_Subtraction(BitMask,BitMask).left.parameter.Out.0\;
                            \BitMask::op_Subtraction(BitMask,BitMask).0.right.parameter.In\ <= \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::op_Subtraction(BitMask,BitMask).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).BitMask::op_Subtraction(BitMask,UInt32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Subtraction(BitMask,BitMask).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).BitMask::op_Subtraction(BitMask,UInt32).0.runningState.0\ := AfterFinished;
                                    \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::op_Subtraction(BitMask,BitMask)._Finished.0\ <= true;
                                    \BitMask::op_Subtraction(BitMask,BitMask).0._Started\ <= false;
                                    \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::op_Subtraction(BitMask,BitMask).return.0\ <= \BitMask::op_Subtraction(BitMask,BitMask).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).BitMask::op_Subtraction(BitMask,UInt32).0.runningState.0\ := WaitingForStarted;
                            \BitMask::op_Subtraction(BitMask,UInt32).0.BitMask::op_Subtraction(BitMask,BitMask)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::AddAlignedFractions(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean).0
                case \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\) then 
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningIndex.0\ := 0;
                            \BitMask::op_Subtraction(BitMask,BitMask).0._Started\ <= true;
                            \BitMask::op_Subtraction(BitMask,BitMask).0.left.parameter.In\ <= \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask).left.parameter.Out.0\;
                            \BitMask::op_Subtraction(BitMask,BitMask).0.right.parameter.In\ <= \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Subtraction(BitMask,BitMask).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningState.0\ := AfterFinished;
                                    \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask)._Finished.0\ <= true;
                                    \BitMask::op_Subtraction(BitMask,BitMask).0._Started\ <= false;
                                    \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask).return.0\ <= \BitMask::op_Subtraction(BitMask,BitMask).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningState.0\ := WaitingForStarted;
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_Subtraction(BitMask,BitMask)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Void Lombiq.Unum.UnumEnvironment::.ctor(System.Byte,System.Byte).0
                case \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\ := 0;
                            \BitMask::op_Subtraction(BitMask,BitMask).0._Started\ <= true;
                            \BitMask::op_Subtraction(BitMask,BitMask).0.left.parameter.In\ <= \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask).left.parameter.Out.0\;
                            \BitMask::op_Subtraction(BitMask,BitMask).0.right.parameter.In\ <= \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Subtraction(BitMask,BitMask).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := AfterFinished;
                                    \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Finished.0\ <= true;
                                    \BitMask::op_Subtraction(BitMask,BitMask).0._Started\ <= false;
                                    \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask).return.0\ <= \BitMask::op_Subtraction(BitMask,BitMask).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,BitMask).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := WaitingForStarted;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,BitMask)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean) start
    \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).BitMask::op_BitwiseOr(BitMask,BitMask).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).BitMask::op_BitwiseOr(BitMask,BitMask).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).BitMask::op_BitwiseAnd(BitMask,BitMask).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).BitMask::op_BitwiseAnd(BitMask,BitMask).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::.ctor(UnumEnvironment).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::.ctor(UnumEnvironment).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::AddExactUnums(Unum,Unum).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).BitMask::op_BitwiseOr(BitMask,BitMask).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).BitMask::op_BitwiseOr(BitMask,BitMask).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).BitMask::op_BitwiseAnd(BitMask,BitMask).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).BitMask::op_BitwiseAnd(BitMask,BitMask).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::.ctor(UnumEnvironment).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::.ctor(UnumEnvironment).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := WaitingForStarted;
                \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= false;
                \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= false;
                \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= false;
                \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= false;
                \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseOr(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0
                case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).BitMask::op_BitwiseOr(BitMask,BitMask).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Started.0\) then 
                            \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).BitMask::op_BitwiseOr(BitMask,BitMask).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).BitMask::op_BitwiseOr(BitMask,BitMask).0.runningIndex.0\ := 0;
                            \BitMask::.ctor(UInt16,Boolean).0._Started\ <= true;
                            \BitMask::.ctor(UInt16,Boolean).0.this.parameter.In\ <= \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\;
                            \BitMask::.ctor(UInt16,Boolean).0.size.parameter.In\ <= \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\;
                            \BitMask::.ctor(UInt16,Boolean).0.allOne.parameter.In\ <= \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).BitMask::op_BitwiseOr(BitMask,BitMask).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::.ctor(UInt16,Boolean).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).BitMask::op_BitwiseOr(BitMask,BitMask).0.runningState.0\ := AfterFinished;
                                    \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= true;
                                    \BitMask::.ctor(UInt16,Boolean).0._Started\ <= false;
                                    \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\ <= \BitMask::.ctor(UInt16,Boolean).0.this.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).BitMask::op_BitwiseOr(BitMask,BitMask).0.runningState.0\ := WaitingForStarted;
                            \BitMask::op_BitwiseOr(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseAnd(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask).0
                case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).BitMask::op_BitwiseAnd(BitMask,BitMask).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Started.0\) then 
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).BitMask::op_BitwiseAnd(BitMask,BitMask).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).BitMask::op_BitwiseAnd(BitMask,BitMask).0.runningIndex.0\ := 0;
                            \BitMask::.ctor(UInt16,Boolean).0._Started\ <= true;
                            \BitMask::.ctor(UInt16,Boolean).0.this.parameter.In\ <= \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\;
                            \BitMask::.ctor(UInt16,Boolean).0.size.parameter.In\ <= \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\;
                            \BitMask::.ctor(UInt16,Boolean).0.allOne.parameter.In\ <= \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).BitMask::op_BitwiseAnd(BitMask,BitMask).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::.ctor(UInt16,Boolean).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).BitMask::op_BitwiseAnd(BitMask,BitMask).0.runningState.0\ := AfterFinished;
                                    \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= true;
                                    \BitMask::.ctor(UInt16,Boolean).0._Started\ <= false;
                                    \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\ <= \BitMask::.ctor(UInt16,Boolean).0.this.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).BitMask::op_BitwiseAnd(BitMask,BitMask).0.runningState.0\ := WaitingForStarted;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment).0
                case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::.ctor(UnumEnvironment).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean)._Started.0\) then 
                            \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::.ctor(UnumEnvironment).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::.ctor(UnumEnvironment).0.runningIndex.0\ := 0;
                            \BitMask::.ctor(UInt16,Boolean).0._Started\ <= true;
                            \BitMask::.ctor(UInt16,Boolean).0.this.parameter.In\ <= \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\;
                            \BitMask::.ctor(UInt16,Boolean).0.size.parameter.In\ <= \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\;
                            \BitMask::.ctor(UInt16,Boolean).0.allOne.parameter.In\ <= \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::.ctor(UnumEnvironment).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::.ctor(UInt16,Boolean).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::.ctor(UnumEnvironment).0.runningState.0\ := AfterFinished;
                                    \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= true;
                                    \BitMask::.ctor(UInt16,Boolean).0._Started\ <= false;
                                    \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\ <= \BitMask::.ctor(UInt16,Boolean).0.this.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::.ctor(UnumEnvironment).0.runningState.0\ := WaitingForStarted;
                            \Unum::.ctor(UnumEnvironment).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0
                case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean)._Started.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                            \BitMask::.ctor(UInt16,Boolean).0._Started\ <= true;
                            \BitMask::.ctor(UInt16,Boolean).0.this.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\;
                            \BitMask::.ctor(UInt16,Boolean).0.size.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\;
                            \BitMask::.ctor(UInt16,Boolean).0.allOne.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::.ctor(UInt16,Boolean).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := AfterFinished;
                                    \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= true;
                                    \BitMask::.ctor(UInt16,Boolean).0._Started\ <= false;
                                    \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\ <= \BitMask::.ctor(UInt16,Boolean).0.this.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::AddAlignedFractions(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean).0
                case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean)._Started.0\) then 
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningIndex.0\ := 0;
                            \BitMask::.ctor(UInt16,Boolean).0._Started\ <= true;
                            \BitMask::.ctor(UInt16,Boolean).0.this.parameter.In\ <= \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\;
                            \BitMask::.ctor(UInt16,Boolean).0.size.parameter.In\ <= \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\;
                            \BitMask::.ctor(UInt16,Boolean).0.allOne.parameter.In\ <= \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::.ctor(UInt16,Boolean).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningState.0\ := AfterFinished;
                                    \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= true;
                                    \BitMask::.ctor(UInt16,Boolean).0._Started\ <= false;
                                    \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\ <= \BitMask::.ctor(UInt16,Boolean).0.this.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.runningState.0\ := WaitingForStarted;
                            \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Void Lombiq.Unum.UnumEnvironment::.ctor(System.Byte,System.Byte).0
                case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\ := 0;
                            \BitMask::.ctor(UInt16,Boolean).0._Started\ <= true;
                            \BitMask::.ctor(UInt16,Boolean).0.this.parameter.In\ <= \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).this.parameter.Out.0\;
                            \BitMask::.ctor(UInt16,Boolean).0.size.parameter.In\ <= \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).size.parameter.Out.0\;
                            \BitMask::.ctor(UInt16,Boolean).0.allOne.parameter.In\ <= \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).allOne.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::.ctor(UInt16,Boolean).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := AfterFinished;
                                    \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= true;
                                    \BitMask::.ctor(UInt16,Boolean).0._Started\ <= false;
                                    \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean).this.parameter.In.0\ <= \BitMask::.ctor(UInt16,Boolean).0.this.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::.ctor(UInt16,Boolean).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := WaitingForStarted;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::.ctor(UInt16,Boolean)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.Void Lombiq.Unum.BitMask::.ctor(System.UInt16,System.Boolean) end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32) start
    \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).BitMask::op_RightShift(BitMask,Int32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).BitMask::op_RightShift(BitMask,Int32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::FractionToUintArray().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::FractionToUintArray().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::FractionMask().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::FractionMask().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::ExponentMask().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::ExponentMask().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::AddExactUnums(Unum,Unum).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).BitMask::op_RightShift(BitMask,Int32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).BitMask::op_RightShift(BitMask,Int32).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::FractionToUintArray().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::FractionToUintArray().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::FractionMask().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::FractionMask().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::ExponentMask().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::ExponentMask().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                \BitMask::op_RightShift(BitMask,Int32).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= false;
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= false;
                \Unum::FractionToUintArray().0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= false;
                \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= false;
                \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_RightShift(Lombiq.Unum.BitMask,System.Int32).0
                case \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).BitMask::op_RightShift(BitMask,Int32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\BitMask::op_RightShift(BitMask,Int32).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\) then 
                            \BitMask::op_RightShift(BitMask,Int32).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).BitMask::op_RightShift(BitMask,Int32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).BitMask::op_RightShift(BitMask,Int32).0.runningIndex.0\ := 0;
                            \BitMask::op_LeftShift(BitMask,Int32).0._Started\ <= true;
                            \BitMask::op_LeftShift(BitMask,Int32).0.left.parameter.In\ <= \BitMask::op_RightShift(BitMask,Int32).0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\;
                            \BitMask::op_LeftShift(BitMask,Int32).0.right.parameter.In\ <= \BitMask::op_RightShift(BitMask,Int32).0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).BitMask::op_RightShift(BitMask,Int32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_LeftShift(BitMask,Int32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).BitMask::op_RightShift(BitMask,Int32).0.runningState.0\ := AfterFinished;
                                    \BitMask::op_RightShift(BitMask,Int32).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= true;
                                    \BitMask::op_LeftShift(BitMask,Int32).0._Started\ <= false;
                                    \BitMask::op_RightShift(BitMask,Int32).0.BitMask::op_LeftShift(BitMask,Int32).return.0\ <= \BitMask::op_LeftShift(BitMask,Int32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\BitMask::op_RightShift(BitMask,Int32).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).BitMask::op_RightShift(BitMask,Int32).0.runningState.0\ := WaitingForStarted;
                            \BitMask::op_RightShift(BitMask,Int32).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::SetUnumBits(System.Boolean,Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean,System.Byte,System.UInt16).0
                case \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\) then 
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\ := 0;
                            \BitMask::op_LeftShift(BitMask,Int32).0._Started\ <= true;
                            \BitMask::op_LeftShift(BitMask,Int32).0.left.parameter.In\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\;
                            \BitMask::op_LeftShift(BitMask,Int32).0.right.parameter.In\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_LeftShift(BitMask,Int32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := AfterFinished;
                                    \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= true;
                                    \BitMask::op_LeftShift(BitMask,Int32).0._Started\ <= false;
                                    \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32).return.0\ <= \BitMask::op_LeftShift(BitMask,Int32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := WaitingForStarted;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.UInt32[] Lombiq.Unum.Unum::FractionToUintArray().0
                case \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::FractionToUintArray().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::FractionToUintArray().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\) then 
                            \Unum::FractionToUintArray().0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::FractionToUintArray().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::FractionToUintArray().0.runningIndex.0\ := 0;
                            \BitMask::op_LeftShift(BitMask,Int32).0._Started\ <= true;
                            \BitMask::op_LeftShift(BitMask,Int32).0.left.parameter.In\ <= \Unum::FractionToUintArray().0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\;
                            \BitMask::op_LeftShift(BitMask,Int32).0.right.parameter.In\ <= \Unum::FractionToUintArray().0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::FractionToUintArray().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_LeftShift(BitMask,Int32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::FractionToUintArray().0.runningState.0\ := AfterFinished;
                                    \Unum::FractionToUintArray().0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= true;
                                    \BitMask::op_LeftShift(BitMask,Int32).0._Started\ <= false;
                                    \Unum::FractionToUintArray().0.BitMask::op_LeftShift(BitMask,Int32).return.0\ <= \BitMask::op_LeftShift(BitMask,Int32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::FractionToUintArray().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::FractionToUintArray().0.runningState.0\ := WaitingForStarted;
                            \Unum::FractionToUintArray().0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionMask().0
                case \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::FractionMask().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\) then 
                            \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::FractionMask().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::FractionMask().0.runningIndex.0\ := 0;
                            \BitMask::op_LeftShift(BitMask,Int32).0._Started\ <= true;
                            \BitMask::op_LeftShift(BitMask,Int32).0.left.parameter.In\ <= \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\;
                            \BitMask::op_LeftShift(BitMask,Int32).0.right.parameter.In\ <= \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::FractionMask().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_LeftShift(BitMask,Int32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::FractionMask().0.runningState.0\ := AfterFinished;
                                    \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= true;
                                    \BitMask::op_LeftShift(BitMask,Int32).0._Started\ <= false;
                                    \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32).return.0\ <= \BitMask::op_LeftShift(BitMask,Int32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::FractionMask().0.runningState.0\ := WaitingForStarted;
                            \Unum::FractionMask().0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentMask().0
                case \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::ExponentMask().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\) then 
                            \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::ExponentMask().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::ExponentMask().0.runningIndex.0\ := 0;
                            \BitMask::op_LeftShift(BitMask,Int32).0._Started\ <= true;
                            \BitMask::op_LeftShift(BitMask,Int32).0.left.parameter.In\ <= \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\;
                            \BitMask::op_LeftShift(BitMask,Int32).0.right.parameter.In\ <= \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::ExponentMask().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_LeftShift(BitMask,Int32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::ExponentMask().0.runningState.0\ := AfterFinished;
                                    \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= true;
                                    \BitMask::op_LeftShift(BitMask,Int32).0._Started\ <= false;
                                    \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32).return.0\ <= \BitMask::op_LeftShift(BitMask,Int32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::ExponentMask().0.runningState.0\ := WaitingForStarted;
                            \Unum::ExponentMask().0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0
                case \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                            \BitMask::op_LeftShift(BitMask,Int32).0._Started\ <= true;
                            \BitMask::op_LeftShift(BitMask,Int32).0.left.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).left.parameter.Out.0\;
                            \BitMask::op_LeftShift(BitMask,Int32).0.right.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_LeftShift(BitMask,Int32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := AfterFinished;
                                    \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= true;
                                    \BitMask::op_LeftShift(BitMask,Int32).0._Started\ <= false;
                                    \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32).return.0\ <= \BitMask::op_LeftShift(BitMask,Int32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_LeftShift(BitMask,Int32).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_LeftShift(BitMask,Int32)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_LeftShift(Lombiq.Unum.BitMask,System.Int32) end


    -- System.Void Hast::InternalInvocationProxy().System.Boolean Lombiq.Unum.BitMask::op_Equality(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask) start
    \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsExact().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsExact().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsPositive().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsPositive().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsNan().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsNan().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsPositiveInfinity().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsPositiveInfinity().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsNegativeInfinity().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsNegativeInfinity().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsExact().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsExact().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsPositive().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsPositive().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsNan().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsNan().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsPositiveInfinity().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsPositiveInfinity().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsNegativeInfinity().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsNegativeInfinity().0.runningState.0\ := WaitingForStarted;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= false;
                \Unum::IsExact().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= false;
                \Unum::IsPositive().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= false;
                \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= false;
                \Unum::IsPositiveInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= false;
                \Unum::IsNegativeInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.UInt32[],System.Boolean).0
                case \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Equality(BitMask,BitMask)._Started.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ := 0;
                            \BitMask::op_Equality(BitMask,BitMask).0._Started\ <= true;
                            \BitMask::op_Equality(BitMask,BitMask).0.left.parameter.In\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Equality(BitMask,BitMask).left.parameter.Out.0\;
                            \BitMask::op_Equality(BitMask,BitMask).0.right.parameter.In\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Equality(BitMask,BitMask).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Equality(BitMask,BitMask).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := AfterFinished;
                                    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= true;
                                    \BitMask::op_Equality(BitMask,BitMask).0._Started\ <= false;
                                    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Equality(BitMask,BitMask).return.0\ <= \BitMask::op_Equality(BitMask,BitMask).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForStarted;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Boolean Lombiq.Unum.Unum::IsExact().0
                case \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsExact().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::IsExact().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\) then 
                            \Unum::IsExact().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsExact().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsExact().0.runningIndex.0\ := 0;
                            \BitMask::op_Equality(BitMask,BitMask).0._Started\ <= true;
                            \BitMask::op_Equality(BitMask,BitMask).0.left.parameter.In\ <= \Unum::IsExact().0.BitMask::op_Equality(BitMask,BitMask).left.parameter.Out.0\;
                            \BitMask::op_Equality(BitMask,BitMask).0.right.parameter.In\ <= \Unum::IsExact().0.BitMask::op_Equality(BitMask,BitMask).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsExact().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Equality(BitMask,BitMask).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsExact().0.runningState.0\ := AfterFinished;
                                    \Unum::IsExact().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= true;
                                    \BitMask::op_Equality(BitMask,BitMask).0._Started\ <= false;
                                    \Unum::IsExact().0.BitMask::op_Equality(BitMask,BitMask).return.0\ <= \BitMask::op_Equality(BitMask,BitMask).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::IsExact().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsExact().0.runningState.0\ := WaitingForStarted;
                            \Unum::IsExact().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Boolean Lombiq.Unum.Unum::IsPositive().0
                case \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsPositive().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::IsPositive().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\) then 
                            \Unum::IsPositive().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsPositive().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsPositive().0.runningIndex.0\ := 0;
                            \BitMask::op_Equality(BitMask,BitMask).0._Started\ <= true;
                            \BitMask::op_Equality(BitMask,BitMask).0.left.parameter.In\ <= \Unum::IsPositive().0.BitMask::op_Equality(BitMask,BitMask).left.parameter.Out.0\;
                            \BitMask::op_Equality(BitMask,BitMask).0.right.parameter.In\ <= \Unum::IsPositive().0.BitMask::op_Equality(BitMask,BitMask).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsPositive().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Equality(BitMask,BitMask).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsPositive().0.runningState.0\ := AfterFinished;
                                    \Unum::IsPositive().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= true;
                                    \BitMask::op_Equality(BitMask,BitMask).0._Started\ <= false;
                                    \Unum::IsPositive().0.BitMask::op_Equality(BitMask,BitMask).return.0\ <= \BitMask::op_Equality(BitMask,BitMask).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::IsPositive().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsPositive().0.runningState.0\ := WaitingForStarted;
                            \Unum::IsPositive().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Boolean Lombiq.Unum.Unum::IsNan().0
                case \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsNan().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\) then 
                            \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsNan().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsNan().0.runningIndex.0\ := 0;
                            \BitMask::op_Equality(BitMask,BitMask).0._Started\ <= true;
                            \BitMask::op_Equality(BitMask,BitMask).0.left.parameter.In\ <= \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask).left.parameter.Out.0\;
                            \BitMask::op_Equality(BitMask,BitMask).0.right.parameter.In\ <= \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsNan().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Equality(BitMask,BitMask).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsNan().0.runningState.0\ := AfterFinished;
                                    \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= true;
                                    \BitMask::op_Equality(BitMask,BitMask).0._Started\ <= false;
                                    \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask).return.0\ <= \BitMask::op_Equality(BitMask,BitMask).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsNan().0.runningState.0\ := WaitingForStarted;
                            \Unum::IsNan().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Boolean Lombiq.Unum.Unum::IsPositiveInfinity().0
                case \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsPositiveInfinity().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::IsPositiveInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\) then 
                            \Unum::IsPositiveInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsPositiveInfinity().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsPositiveInfinity().0.runningIndex.0\ := 0;
                            \BitMask::op_Equality(BitMask,BitMask).0._Started\ <= true;
                            \BitMask::op_Equality(BitMask,BitMask).0.left.parameter.In\ <= \Unum::IsPositiveInfinity().0.BitMask::op_Equality(BitMask,BitMask).left.parameter.Out.0\;
                            \BitMask::op_Equality(BitMask,BitMask).0.right.parameter.In\ <= \Unum::IsPositiveInfinity().0.BitMask::op_Equality(BitMask,BitMask).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsPositiveInfinity().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Equality(BitMask,BitMask).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsPositiveInfinity().0.runningState.0\ := AfterFinished;
                                    \Unum::IsPositiveInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= true;
                                    \BitMask::op_Equality(BitMask,BitMask).0._Started\ <= false;
                                    \Unum::IsPositiveInfinity().0.BitMask::op_Equality(BitMask,BitMask).return.0\ <= \BitMask::op_Equality(BitMask,BitMask).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::IsPositiveInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsPositiveInfinity().0.runningState.0\ := WaitingForStarted;
                            \Unum::IsPositiveInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Boolean Lombiq.Unum.Unum::IsNegativeInfinity().0
                case \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsNegativeInfinity().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::IsNegativeInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\) then 
                            \Unum::IsNegativeInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsNegativeInfinity().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsNegativeInfinity().0.runningIndex.0\ := 0;
                            \BitMask::op_Equality(BitMask,BitMask).0._Started\ <= true;
                            \BitMask::op_Equality(BitMask,BitMask).0.left.parameter.In\ <= \Unum::IsNegativeInfinity().0.BitMask::op_Equality(BitMask,BitMask).left.parameter.Out.0\;
                            \BitMask::op_Equality(BitMask,BitMask).0.right.parameter.In\ <= \Unum::IsNegativeInfinity().0.BitMask::op_Equality(BitMask,BitMask).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsNegativeInfinity().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Equality(BitMask,BitMask).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsNegativeInfinity().0.runningState.0\ := AfterFinished;
                                    \Unum::IsNegativeInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= true;
                                    \BitMask::op_Equality(BitMask,BitMask).0._Started\ <= false;
                                    \Unum::IsNegativeInfinity().0.BitMask::op_Equality(BitMask,BitMask).return.0\ <= \BitMask::op_Equality(BitMask,BitMask).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::IsNegativeInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Equality(BitMask,BitMask).Unum::IsNegativeInfinity().0.runningState.0\ := WaitingForStarted;
                            \Unum::IsNegativeInfinity().0.BitMask::op_Equality(BitMask,BitMask)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.Boolean Lombiq.Unum.BitMask::op_Equality(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask) end


    -- System.Void Hast::InternalInvocationProxy().System.UInt16 Lombiq.Unum.Unum::get_Size() start
    \Hast::InternalInvocationProxy().Unum::get_Size()\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Unum::get_Size().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::get_Size().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Unum::get_Size().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::get_Size().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Unum::get_Size().Unum::FractionMask().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::get_Size().Unum::FractionMask().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Unum::get_Size().Unum::ExponentMask().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::get_Size().Unum::ExponentMask().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Unum::get_Size().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::get_Size().Unum::AddExactUnums(Unum,Unum).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().Unum::get_Size().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::get_Size().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Unum::get_Size().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::get_Size().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Unum::get_Size().Unum::FractionMask().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::get_Size().Unum::FractionMask().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Unum::get_Size().Unum::ExponentMask().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::get_Size().Unum::ExponentMask().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Unum::get_Size().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::get_Size().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size()._Finished.0\ <= false;
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_Size()._Finished.0\ <= false;
                \Unum::FractionMask().0.Unum::get_Size()._Finished.0\ <= false;
                \Unum::ExponentMask().0.Unum::get_Size()._Finished.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::get_Size()._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.UInt32[],System.Boolean).0
                case \Hast::InternalInvocationProxy().Unum::get_Size().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size()._Started.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::get_Size().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::get_Size().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ := 0;
                            \Unum::get_Size().0._Started\ <= true;
                            \Unum::get_Size().0.this.parameter.In\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::get_Size().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::get_Size().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::get_Size().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := AfterFinished;
                                    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size()._Finished.0\ <= true;
                                    \Unum::get_Size().0._Started\ <= false;
                                    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size().return.0\ <= \Unum::get_Size().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::get_Size().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForStarted;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::get_Size()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::SetUnumBits(System.Boolean,Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean,System.Byte,System.UInt16).0
                case \Hast::InternalInvocationProxy().Unum::get_Size().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_Size()._Started.0\) then 
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_Size()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::get_Size().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::get_Size().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\ := 0;
                            \Unum::get_Size().0._Started\ <= true;
                            \Unum::get_Size().0.this.parameter.In\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_Size().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::get_Size().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::get_Size().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::get_Size().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := AfterFinished;
                                    \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_Size()._Finished.0\ <= true;
                                    \Unum::get_Size().0._Started\ <= false;
                                    \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_Size().return.0\ <= \Unum::get_Size().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_Size()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::get_Size().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := WaitingForStarted;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_Size()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionMask().0
                case \Hast::InternalInvocationProxy().Unum::get_Size().Unum::FractionMask().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::FractionMask().0.Unum::get_Size()._Started.0\) then 
                            \Unum::FractionMask().0.Unum::get_Size()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::get_Size().Unum::FractionMask().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::get_Size().Unum::FractionMask().0.runningIndex.0\ := 0;
                            \Unum::get_Size().0._Started\ <= true;
                            \Unum::get_Size().0.this.parameter.In\ <= \Unum::FractionMask().0.Unum::get_Size().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::get_Size().Unum::FractionMask().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::get_Size().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::get_Size().Unum::FractionMask().0.runningState.0\ := AfterFinished;
                                    \Unum::FractionMask().0.Unum::get_Size()._Finished.0\ <= true;
                                    \Unum::get_Size().0._Started\ <= false;
                                    \Unum::FractionMask().0.Unum::get_Size().return.0\ <= \Unum::get_Size().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::FractionMask().0.Unum::get_Size()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::get_Size().Unum::FractionMask().0.runningState.0\ := WaitingForStarted;
                            \Unum::FractionMask().0.Unum::get_Size()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentMask().0
                case \Hast::InternalInvocationProxy().Unum::get_Size().Unum::ExponentMask().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::ExponentMask().0.Unum::get_Size()._Started.0\) then 
                            \Unum::ExponentMask().0.Unum::get_Size()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::get_Size().Unum::ExponentMask().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::get_Size().Unum::ExponentMask().0.runningIndex.0\ := 0;
                            \Unum::get_Size().0._Started\ <= true;
                            \Unum::get_Size().0.this.parameter.In\ <= \Unum::ExponentMask().0.Unum::get_Size().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::get_Size().Unum::ExponentMask().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::get_Size().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::get_Size().Unum::ExponentMask().0.runningState.0\ := AfterFinished;
                                    \Unum::ExponentMask().0.Unum::get_Size()._Finished.0\ <= true;
                                    \Unum::get_Size().0._Started\ <= false;
                                    \Unum::ExponentMask().0.Unum::get_Size().return.0\ <= \Unum::get_Size().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::ExponentMask().0.Unum::get_Size()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::get_Size().Unum::ExponentMask().0.runningState.0\ := WaitingForStarted;
                            \Unum::ExponentMask().0.Unum::get_Size()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0
                case \Hast::InternalInvocationProxy().Unum::get_Size().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::get_Size()._Started.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_Size()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::get_Size().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::get_Size().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                            \Unum::get_Size().0._Started\ <= true;
                            \Unum::get_Size().0.this.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::get_Size().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::get_Size().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::get_Size().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::get_Size().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := AfterFinished;
                                    \Unum::AddExactUnums(Unum,Unum).0.Unum::get_Size()._Finished.0\ <= true;
                                    \Unum::get_Size().0._Started\ <= false;
                                    \Unum::AddExactUnums(Unum,Unum).0.Unum::get_Size().return.0\ <= \Unum::get_Size().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::get_Size()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::get_Size().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_Size()._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.UInt16 Lombiq.Unum.Unum::get_Size() end


    -- System.Void Hast::InternalInvocationProxy().System.UInt16 Lombiq.Unum.BitMask::GetMostSignificantOnePosition() start
    \Hast::InternalInvocationProxy().BitMask::GetMostSignificantOnePosition()\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().BitMask::GetMostSignificantOnePosition().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::GetMostSignificantOnePosition().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::GetMostSignificantOnePosition().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::GetMostSignificantOnePosition().Unum::AddExactUnums(Unum,Unum).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().BitMask::GetMostSignificantOnePosition().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::GetMostSignificantOnePosition().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::GetMostSignificantOnePosition().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::GetMostSignificantOnePosition().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition()._Finished.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.UInt32[],System.Boolean).0
                case \Hast::InternalInvocationProxy().BitMask::GetMostSignificantOnePosition().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition()._Started.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::GetMostSignificantOnePosition().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::GetMostSignificantOnePosition().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ := 0;
                            \BitMask::GetMostSignificantOnePosition().0._Started\ <= true;
                            \BitMask::GetMostSignificantOnePosition().0.this.parameter.In\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::GetMostSignificantOnePosition().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::GetMostSignificantOnePosition().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::GetMostSignificantOnePosition().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := AfterFinished;
                                    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition()._Finished.0\ <= true;
                                    \BitMask::GetMostSignificantOnePosition().0._Started\ <= false;
                                    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition().return.0\ <= \BitMask::GetMostSignificantOnePosition().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::GetMostSignificantOnePosition().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForStarted;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetMostSignificantOnePosition()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0
                case \Hast::InternalInvocationProxy().BitMask::GetMostSignificantOnePosition().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Started.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::GetMostSignificantOnePosition().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::GetMostSignificantOnePosition().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                            \BitMask::GetMostSignificantOnePosition().0._Started\ <= true;
                            \BitMask::GetMostSignificantOnePosition().0.this.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::GetMostSignificantOnePosition().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::GetMostSignificantOnePosition().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::GetMostSignificantOnePosition().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := AfterFinished;
                                    \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Finished.0\ <= true;
                                    \BitMask::GetMostSignificantOnePosition().0._Started\ <= false;
                                    \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition().return.0\ <= \BitMask::GetMostSignificantOnePosition().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::GetMostSignificantOnePosition().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::GetMostSignificantOnePosition()._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.UInt16 Lombiq.Unum.BitMask::GetMostSignificantOnePosition() end


    -- System.Void Hast::InternalInvocationProxy().System.UInt32 Lombiq.Unum.BitMask::GetLowest32Bits() start
    \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits()\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::ExponentSize().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::ExponentSize().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::FractionSize().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::FractionSize().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::HiddenBitIsOne().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::HiddenBitIsOne().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::ExponentValueWithBias().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::ExponentValueWithBias().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::ExponentSize().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::ExponentSize().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::FractionSize().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::FractionSize().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::HiddenBitIsOne().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::HiddenBitIsOne().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::ExponentValueWithBias().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::ExponentValueWithBias().0.runningState.0\ := WaitingForStarted;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits()._Finished.0\ <= false;
                \Unum::ExponentSize().0.BitMask::GetLowest32Bits()._Finished.0\ <= false;
                \Unum::FractionSize().0.BitMask::GetLowest32Bits()._Finished.0\ <= false;
                \Unum::HiddenBitIsOne().0.BitMask::GetLowest32Bits()._Finished.0\ <= false;
                \Unum::ExponentValueWithBias().0.BitMask::GetLowest32Bits()._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.UInt32[],System.Boolean).0
                case \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits()._Started.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ := 0;
                            \BitMask::GetLowest32Bits().0._Started\ <= true;
                            \BitMask::GetLowest32Bits().0.this.parameter.In\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::GetLowest32Bits().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := AfterFinished;
                                    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits()._Finished.0\ <= true;
                                    \BitMask::GetLowest32Bits().0._Started\ <= false;
                                    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits().return.0\ <= \BitMask::GetLowest32Bits().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForStarted;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::GetLowest32Bits()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Byte Lombiq.Unum.Unum::ExponentSize().0
                case \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::ExponentSize().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::ExponentSize().0.BitMask::GetLowest32Bits()._Started.0\) then 
                            \Unum::ExponentSize().0.BitMask::GetLowest32Bits()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::ExponentSize().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::ExponentSize().0.runningIndex.0\ := 0;
                            \BitMask::GetLowest32Bits().0._Started\ <= true;
                            \BitMask::GetLowest32Bits().0.this.parameter.In\ <= \Unum::ExponentSize().0.BitMask::GetLowest32Bits().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::ExponentSize().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::GetLowest32Bits().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::ExponentSize().0.runningState.0\ := AfterFinished;
                                    \Unum::ExponentSize().0.BitMask::GetLowest32Bits()._Finished.0\ <= true;
                                    \BitMask::GetLowest32Bits().0._Started\ <= false;
                                    \Unum::ExponentSize().0.BitMask::GetLowest32Bits().return.0\ <= \BitMask::GetLowest32Bits().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::ExponentSize().0.BitMask::GetLowest32Bits()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::ExponentSize().0.runningState.0\ := WaitingForStarted;
                            \Unum::ExponentSize().0.BitMask::GetLowest32Bits()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.UInt16 Lombiq.Unum.Unum::FractionSize().0
                case \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::FractionSize().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::FractionSize().0.BitMask::GetLowest32Bits()._Started.0\) then 
                            \Unum::FractionSize().0.BitMask::GetLowest32Bits()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::FractionSize().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::FractionSize().0.runningIndex.0\ := 0;
                            \BitMask::GetLowest32Bits().0._Started\ <= true;
                            \BitMask::GetLowest32Bits().0.this.parameter.In\ <= \Unum::FractionSize().0.BitMask::GetLowest32Bits().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::FractionSize().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::GetLowest32Bits().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::FractionSize().0.runningState.0\ := AfterFinished;
                                    \Unum::FractionSize().0.BitMask::GetLowest32Bits()._Finished.0\ <= true;
                                    \BitMask::GetLowest32Bits().0._Started\ <= false;
                                    \Unum::FractionSize().0.BitMask::GetLowest32Bits().return.0\ <= \BitMask::GetLowest32Bits().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::FractionSize().0.BitMask::GetLowest32Bits()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::FractionSize().0.runningState.0\ := WaitingForStarted;
                            \Unum::FractionSize().0.BitMask::GetLowest32Bits()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Boolean Lombiq.Unum.Unum::HiddenBitIsOne().0
                case \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::HiddenBitIsOne().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::HiddenBitIsOne().0.BitMask::GetLowest32Bits()._Started.0\) then 
                            \Unum::HiddenBitIsOne().0.BitMask::GetLowest32Bits()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::HiddenBitIsOne().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::HiddenBitIsOne().0.runningIndex.0\ := 0;
                            \BitMask::GetLowest32Bits().0._Started\ <= true;
                            \BitMask::GetLowest32Bits().0.this.parameter.In\ <= \Unum::HiddenBitIsOne().0.BitMask::GetLowest32Bits().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::HiddenBitIsOne().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::GetLowest32Bits().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::HiddenBitIsOne().0.runningState.0\ := AfterFinished;
                                    \Unum::HiddenBitIsOne().0.BitMask::GetLowest32Bits()._Finished.0\ <= true;
                                    \BitMask::GetLowest32Bits().0._Started\ <= false;
                                    \Unum::HiddenBitIsOne().0.BitMask::GetLowest32Bits().return.0\ <= \BitMask::GetLowest32Bits().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::HiddenBitIsOne().0.BitMask::GetLowest32Bits()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::HiddenBitIsOne().0.runningState.0\ := WaitingForStarted;
                            \Unum::HiddenBitIsOne().0.BitMask::GetLowest32Bits()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Int32 Lombiq.Unum.Unum::ExponentValueWithBias().0
                case \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::ExponentValueWithBias().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::ExponentValueWithBias().0.BitMask::GetLowest32Bits()._Started.0\) then 
                            \Unum::ExponentValueWithBias().0.BitMask::GetLowest32Bits()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::ExponentValueWithBias().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::ExponentValueWithBias().0.runningIndex.0\ := 0;
                            \BitMask::GetLowest32Bits().0._Started\ <= true;
                            \BitMask::GetLowest32Bits().0.this.parameter.In\ <= \Unum::ExponentValueWithBias().0.BitMask::GetLowest32Bits().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::ExponentValueWithBias().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::GetLowest32Bits().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::ExponentValueWithBias().0.runningState.0\ := AfterFinished;
                                    \Unum::ExponentValueWithBias().0.BitMask::GetLowest32Bits()._Finished.0\ <= true;
                                    \BitMask::GetLowest32Bits().0._Started\ <= false;
                                    \Unum::ExponentValueWithBias().0.BitMask::GetLowest32Bits().return.0\ <= \BitMask::GetLowest32Bits().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::ExponentValueWithBias().0.BitMask::GetLowest32Bits()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::GetLowest32Bits().Unum::ExponentValueWithBias().0.runningState.0\ := WaitingForStarted;
                            \Unum::ExponentValueWithBias().0.BitMask::GetLowest32Bits()._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.UInt32 Lombiq.Unum.BitMask::GetLowest32Bits() end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,System.UInt32) start
    \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::ExponentSize().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::ExponentSize().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::FractionSize().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::FractionSize().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::ExponentSize().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::ExponentSize().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::FractionSize().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::FractionSize().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := WaitingForStarted;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= false;
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= false;
                \Unum::ExponentSize().0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= false;
                \Unum::FractionSize().0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= false;
                \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= false;
                \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.UInt32[],System.Boolean).0
                case \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ := 0;
                            \BitMask::op_Addition(BitMask,UInt32).0._Started\ <= true;
                            \BitMask::op_Addition(BitMask,UInt32).0.left.parameter.In\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Addition(BitMask,UInt32).left.parameter.Out.0\;
                            \BitMask::op_Addition(BitMask,UInt32).0.right.parameter.In\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Addition(BitMask,UInt32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := AfterFinished;
                                    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= true;
                                    \BitMask::op_Addition(BitMask,UInt32).0._Started\ <= false;
                                    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Addition(BitMask,UInt32).return.0\ <= \BitMask::op_Addition(BitMask,UInt32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForStarted;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::SetUnumBits(System.Boolean,Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean,System.Byte,System.UInt16).0
                case \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\) then 
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\ := 0;
                            \BitMask::op_Addition(BitMask,UInt32).0._Started\ <= true;
                            \BitMask::op_Addition(BitMask,UInt32).0.left.parameter.In\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,UInt32).left.parameter.Out.0\;
                            \BitMask::op_Addition(BitMask,UInt32).0.right.parameter.In\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Addition(BitMask,UInt32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := AfterFinished;
                                    \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= true;
                                    \BitMask::op_Addition(BitMask,UInt32).0._Started\ <= false;
                                    \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,UInt32).return.0\ <= \BitMask::op_Addition(BitMask,UInt32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := WaitingForStarted;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Byte Lombiq.Unum.Unum::ExponentSize().0
                case \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::ExponentSize().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::ExponentSize().0.BitMask::op_Addition(BitMask,UInt32)._Started.0\) then 
                            \Unum::ExponentSize().0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::ExponentSize().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::ExponentSize().0.runningIndex.0\ := 0;
                            \BitMask::op_Addition(BitMask,UInt32).0._Started\ <= true;
                            \BitMask::op_Addition(BitMask,UInt32).0.left.parameter.In\ <= \Unum::ExponentSize().0.BitMask::op_Addition(BitMask,UInt32).left.parameter.Out.0\;
                            \BitMask::op_Addition(BitMask,UInt32).0.right.parameter.In\ <= \Unum::ExponentSize().0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::ExponentSize().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Addition(BitMask,UInt32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::ExponentSize().0.runningState.0\ := AfterFinished;
                                    \Unum::ExponentSize().0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= true;
                                    \BitMask::op_Addition(BitMask,UInt32).0._Started\ <= false;
                                    \Unum::ExponentSize().0.BitMask::op_Addition(BitMask,UInt32).return.0\ <= \BitMask::op_Addition(BitMask,UInt32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::ExponentSize().0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::ExponentSize().0.runningState.0\ := WaitingForStarted;
                            \Unum::ExponentSize().0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.UInt16 Lombiq.Unum.Unum::FractionSize().0
                case \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::FractionSize().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::FractionSize().0.BitMask::op_Addition(BitMask,UInt32)._Started.0\) then 
                            \Unum::FractionSize().0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::FractionSize().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::FractionSize().0.runningIndex.0\ := 0;
                            \BitMask::op_Addition(BitMask,UInt32).0._Started\ <= true;
                            \BitMask::op_Addition(BitMask,UInt32).0.left.parameter.In\ <= \Unum::FractionSize().0.BitMask::op_Addition(BitMask,UInt32).left.parameter.Out.0\;
                            \BitMask::op_Addition(BitMask,UInt32).0.right.parameter.In\ <= \Unum::FractionSize().0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::FractionSize().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Addition(BitMask,UInt32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::FractionSize().0.runningState.0\ := AfterFinished;
                                    \Unum::FractionSize().0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= true;
                                    \BitMask::op_Addition(BitMask,UInt32).0._Started\ <= false;
                                    \Unum::FractionSize().0.BitMask::op_Addition(BitMask,UInt32).return.0\ <= \BitMask::op_Addition(BitMask,UInt32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::FractionSize().0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::FractionSize().0.runningState.0\ := WaitingForStarted;
                            \Unum::FractionSize().0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentValueToExponentBits(System.Int32,System.Byte).0
                case \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\) then 
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningIndex.0\ := 0;
                            \BitMask::op_Addition(BitMask,UInt32).0._Started\ <= true;
                            \BitMask::op_Addition(BitMask,UInt32).0.left.parameter.In\ <= \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32).left.parameter.Out.0\;
                            \BitMask::op_Addition(BitMask,UInt32).0.right.parameter.In\ <= \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Addition(BitMask,UInt32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningState.0\ := AfterFinished;
                                    \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= true;
                                    \BitMask::op_Addition(BitMask,UInt32).0._Started\ <= false;
                                    \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32).return.0\ <= \BitMask::op_Addition(BitMask,UInt32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningState.0\ := WaitingForStarted;
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Void Lombiq.Unum.UnumEnvironment::.ctor(System.Byte,System.Byte).0
                case \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\ := 0;
                            \BitMask::op_Addition(BitMask,UInt32).0._Started\ <= true;
                            \BitMask::op_Addition(BitMask,UInt32).0.left.parameter.In\ <= \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,UInt32).left.parameter.Out.0\;
                            \BitMask::op_Addition(BitMask,UInt32).0.right.parameter.In\ <= \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,UInt32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Addition(BitMask,UInt32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := AfterFinished;
                                    \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= true;
                                    \BitMask::op_Addition(BitMask,UInt32).0._Started\ <= false;
                                    \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,UInt32).return.0\ <= \BitMask::op_Addition(BitMask,UInt32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Addition(BitMask,UInt32).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := WaitingForStarted;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Addition(BitMask,UInt32)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Addition(Lombiq.Unum.BitMask,System.UInt32) end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::ShiftOutLeastSignificantZeros() start
    \Hast::InternalInvocationProxy().BitMask::ShiftOutLeastSignificantZeros()\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().BitMask::ShiftOutLeastSignificantZeros().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::ShiftOutLeastSignificantZeros().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::ShiftOutLeastSignificantZeros().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::ShiftOutLeastSignificantZeros().Unum::AddExactUnums(Unum,Unum).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().BitMask::ShiftOutLeastSignificantZeros().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::ShiftOutLeastSignificantZeros().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::ShiftOutLeastSignificantZeros().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::ShiftOutLeastSignificantZeros().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::ShiftOutLeastSignificantZeros()._Finished.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.BitMask::ShiftOutLeastSignificantZeros()._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.UInt32[],System.Boolean).0
                case \Hast::InternalInvocationProxy().BitMask::ShiftOutLeastSignificantZeros().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::ShiftOutLeastSignificantZeros()._Started.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::ShiftOutLeastSignificantZeros()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::ShiftOutLeastSignificantZeros().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::ShiftOutLeastSignificantZeros().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ := 0;
                            \BitMask::ShiftOutLeastSignificantZeros().0._Started\ <= true;
                            \BitMask::ShiftOutLeastSignificantZeros().0.this.parameter.In\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::ShiftOutLeastSignificantZeros().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::ShiftOutLeastSignificantZeros().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::ShiftOutLeastSignificantZeros().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::ShiftOutLeastSignificantZeros().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := AfterFinished;
                                    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::ShiftOutLeastSignificantZeros()._Finished.0\ <= true;
                                    \BitMask::ShiftOutLeastSignificantZeros().0._Started\ <= false;
                                    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::ShiftOutLeastSignificantZeros().return.0\ <= \BitMask::ShiftOutLeastSignificantZeros().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::ShiftOutLeastSignificantZeros()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::ShiftOutLeastSignificantZeros().Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForStarted;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::ShiftOutLeastSignificantZeros()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0
                case \Hast::InternalInvocationProxy().BitMask::ShiftOutLeastSignificantZeros().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::ShiftOutLeastSignificantZeros()._Started.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::ShiftOutLeastSignificantZeros()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::ShiftOutLeastSignificantZeros().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::ShiftOutLeastSignificantZeros().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                            \BitMask::ShiftOutLeastSignificantZeros().0._Started\ <= true;
                            \BitMask::ShiftOutLeastSignificantZeros().0.this.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.BitMask::ShiftOutLeastSignificantZeros().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::ShiftOutLeastSignificantZeros().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::ShiftOutLeastSignificantZeros().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::ShiftOutLeastSignificantZeros().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := AfterFinished;
                                    \Unum::AddExactUnums(Unum,Unum).0.BitMask::ShiftOutLeastSignificantZeros()._Finished.0\ <= true;
                                    \BitMask::ShiftOutLeastSignificantZeros().0._Started\ <= false;
                                    \Unum::AddExactUnums(Unum,Unum).0.BitMask::ShiftOutLeastSignificantZeros().return.0\ <= \BitMask::ShiftOutLeastSignificantZeros().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::ShiftOutLeastSignificantZeros()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::ShiftOutLeastSignificantZeros().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::ShiftOutLeastSignificantZeros()._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::ShiftOutLeastSignificantZeros() end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetZero(System.UInt16) start
    \Hast::InternalInvocationProxy().BitMask::SetZero(UInt16)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().BitMask::SetZero(UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::SetZero(UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::SetZero(UInt16).Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::SetZero(UInt16).Unum::AddExactUnums(Unum,Unum).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().BitMask::SetZero(UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::SetZero(UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::SetZero(UInt16).Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::SetZero(UInt16).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::SetZero(UInt16)._Finished.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.BitMask::SetZero(UInt16)._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.UInt32[],System.Boolean).0
                case \Hast::InternalInvocationProxy().BitMask::SetZero(UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::SetZero(UInt16)._Started.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::SetZero(UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::SetZero(UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::SetZero(UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ := 0;
                            \BitMask::SetZero(UInt16).0._Started\ <= true;
                            \BitMask::SetZero(UInt16).0.this.parameter.In\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::SetZero(UInt16).this.parameter.Out.0\;
                            \BitMask::SetZero(UInt16).0.index.parameter.In\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::SetZero(UInt16).index.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::SetZero(UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::SetZero(UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::SetZero(UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := AfterFinished;
                                    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::SetZero(UInt16)._Finished.0\ <= true;
                                    \BitMask::SetZero(UInt16).0._Started\ <= false;
                                    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::SetZero(UInt16).return.0\ <= \BitMask::SetZero(UInt16).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::SetZero(UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::SetZero(UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForStarted;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.BitMask::SetZero(UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0
                case \Hast::InternalInvocationProxy().BitMask::SetZero(UInt16).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::SetZero(UInt16)._Started.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::SetZero(UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::SetZero(UInt16).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::SetZero(UInt16).Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                            \BitMask::SetZero(UInt16).0._Started\ <= true;
                            \BitMask::SetZero(UInt16).0.this.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.BitMask::SetZero(UInt16).this.parameter.Out.0\;
                            \BitMask::SetZero(UInt16).0.index.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.BitMask::SetZero(UInt16).index.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::SetZero(UInt16).Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::SetZero(UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::SetZero(UInt16).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := AfterFinished;
                                    \Unum::AddExactUnums(Unum,Unum).0.BitMask::SetZero(UInt16)._Finished.0\ <= true;
                                    \BitMask::SetZero(UInt16).0._Started\ <= false;
                                    \Unum::AddExactUnums(Unum,Unum).0.BitMask::SetZero(UInt16).return.0\ <= \BitMask::SetZero(UInt16).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::AddExactUnums(Unum,Unum).0.BitMask::SetZero(UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::SetZero(UInt16).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                            \Unum::AddExactUnums(Unum,Unum).0.BitMask::SetZero(UInt16)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetZero(System.UInt16) end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::SetUnumBits(System.Boolean,Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean,System.Byte,System.UInt16) start
    \Hast::InternalInvocationProxy().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).Unum::AddExactUnums(Unum,Unum).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Finished.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.UInt32[],System.Boolean).0
                case \Hast::InternalInvocationProxy().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Started.0\) then 
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ := 0;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._Started\ <= true;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.this.parameter.In\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).this.parameter.Out.0\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.signBit.parameter.In\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).signBit.parameter.Out.0\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.exponent.parameter.In\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).exponent.parameter.Out.0\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.fraction.parameter.In\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).fraction.parameter.Out.0\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.uncertainityBit.parameter.In\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).uncertainityBit.parameter.Out.0\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.exponentSize.parameter.In\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).exponentSize.parameter.Out.0\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.fractionSize.parameter.In\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).fractionSize.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := AfterFinished;
                                    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Finished.0\ <= true;
                                    \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._Started\ <= false;
                                    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).return.0\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.runningState.0\ := WaitingForStarted;
                            \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0
                case \Hast::InternalInvocationProxy().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Started.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._Started\ <= true;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.this.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).this.parameter.Out.0\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.signBit.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).signBit.parameter.Out.0\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.exponent.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).exponent.parameter.Out.0\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.fraction.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).fraction.parameter.Out.0\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.uncertainityBit.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).uncertainityBit.parameter.Out.0\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.exponentSize.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).exponentSize.parameter.Out.0\;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.fractionSize.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).fractionSize.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := AfterFinished;
                                    \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Finished.0\ <= true;
                                    \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0._Started\ <= false;
                                    \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).return.0\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::SetUnumBits(System.Boolean,Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean,System.Byte,System.UInt16) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.UInt32[],System.Boolean) start
    -- Signal connections for System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.Int32).0 (#0):
    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._Started\ <= \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean)._Started.0\;
    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.this.parameter.In\ <= \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).this.parameter.Out.0\;
    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.environment.parameter.In\ <= \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).environment.parameter.Out.0\;
    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.value.parameter.In\ <= \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).value.parameter.Out.0\;
    \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.negative.parameter.In\ <= \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).negative.parameter.Out.0\;
    \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean)._Finished.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0._Finished\;
    \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).this.parameter.In.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.this.parameter.Out\;
    \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).environment.parameter.In.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.environment.parameter.Out\;
    \Unum::.ctor(UnumEnvironment,Int32).0.Unum::.ctor(UnumEnvironment,UInt32[],Boolean).value.parameter.In.0\ <= \Unum::.ctor(UnumEnvironment,UInt32[],Boolean).0.value.parameter.Out\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,System.UInt32[],System.Boolean) end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_UncertaintyBitMask() start
    \Hast::InternalInvocationProxy().Unum::get_UncertaintyBitMask()\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Unum::get_UncertaintyBitMask().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::get_UncertaintyBitMask().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Unum::get_UncertaintyBitMask().Unum::IsExact().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::get_UncertaintyBitMask().Unum::IsExact().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().Unum::get_UncertaintyBitMask().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::get_UncertaintyBitMask().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Unum::get_UncertaintyBitMask().Unum::IsExact().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::get_UncertaintyBitMask().Unum::IsExact().0.runningState.0\ := WaitingForStarted;
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_UncertaintyBitMask()._Finished.0\ <= false;
                \Unum::IsExact().0.Unum::get_UncertaintyBitMask()._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::SetUnumBits(System.Boolean,Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean,System.Byte,System.UInt16).0
                case \Hast::InternalInvocationProxy().Unum::get_UncertaintyBitMask().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_UncertaintyBitMask()._Started.0\) then 
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_UncertaintyBitMask()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::get_UncertaintyBitMask().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::get_UncertaintyBitMask().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\ := 0;
                            \Unum::get_UncertaintyBitMask().0._Started\ <= true;
                            \Unum::get_UncertaintyBitMask().0.this.parameter.In\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_UncertaintyBitMask().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::get_UncertaintyBitMask().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::get_UncertaintyBitMask().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::get_UncertaintyBitMask().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := AfterFinished;
                                    \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_UncertaintyBitMask()._Finished.0\ <= true;
                                    \Unum::get_UncertaintyBitMask().0._Started\ <= false;
                                    \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_UncertaintyBitMask().return.0\ <= \Unum::get_UncertaintyBitMask().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_UncertaintyBitMask()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::get_UncertaintyBitMask().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := WaitingForStarted;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_UncertaintyBitMask()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Boolean Lombiq.Unum.Unum::IsExact().0
                case \Hast::InternalInvocationProxy().Unum::get_UncertaintyBitMask().Unum::IsExact().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::IsExact().0.Unum::get_UncertaintyBitMask()._Started.0\) then 
                            \Unum::IsExact().0.Unum::get_UncertaintyBitMask()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::get_UncertaintyBitMask().Unum::IsExact().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::get_UncertaintyBitMask().Unum::IsExact().0.runningIndex.0\ := 0;
                            \Unum::get_UncertaintyBitMask().0._Started\ <= true;
                            \Unum::get_UncertaintyBitMask().0.this.parameter.In\ <= \Unum::IsExact().0.Unum::get_UncertaintyBitMask().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::get_UncertaintyBitMask().Unum::IsExact().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::get_UncertaintyBitMask().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::get_UncertaintyBitMask().Unum::IsExact().0.runningState.0\ := AfterFinished;
                                    \Unum::IsExact().0.Unum::get_UncertaintyBitMask()._Finished.0\ <= true;
                                    \Unum::get_UncertaintyBitMask().0._Started\ <= false;
                                    \Unum::IsExact().0.Unum::get_UncertaintyBitMask().return.0\ <= \Unum::get_UncertaintyBitMask().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::IsExact().0.Unum::get_UncertaintyBitMask()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::get_UncertaintyBitMask().Unum::IsExact().0.runningState.0\ := WaitingForStarted;
                            \Unum::IsExact().0.Unum::get_UncertaintyBitMask()._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_UncertaintyBitMask() end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_SignBitMask() start
    \Hast::InternalInvocationProxy().Unum::get_SignBitMask()\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Unum::get_SignBitMask().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::get_SignBitMask().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Unum::get_SignBitMask().Unum::IsPositive().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::get_SignBitMask().Unum::IsPositive().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().Unum::get_SignBitMask().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::get_SignBitMask().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Unum::get_SignBitMask().Unum::IsPositive().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::get_SignBitMask().Unum::IsPositive().0.runningState.0\ := WaitingForStarted;
                \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_SignBitMask()._Finished.0\ <= false;
                \Unum::IsPositive().0.Unum::get_SignBitMask()._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::SetUnumBits(System.Boolean,Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean,System.Byte,System.UInt16).0
                case \Hast::InternalInvocationProxy().Unum::get_SignBitMask().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_SignBitMask()._Started.0\) then 
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_SignBitMask()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::get_SignBitMask().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::get_SignBitMask().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\ := 0;
                            \Unum::get_SignBitMask().0._Started\ <= true;
                            \Unum::get_SignBitMask().0.this.parameter.In\ <= \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_SignBitMask().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::get_SignBitMask().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::get_SignBitMask().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::get_SignBitMask().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := AfterFinished;
                                    \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_SignBitMask()._Finished.0\ <= true;
                                    \Unum::get_SignBitMask().0._Started\ <= false;
                                    \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_SignBitMask().return.0\ <= \Unum::get_SignBitMask().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_SignBitMask()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::get_SignBitMask().Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.runningState.0\ := WaitingForStarted;
                            \Unum::SetUnumBits(Boolean,BitMask,BitMask,Boolean,Byte,UInt16).0.Unum::get_SignBitMask()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Boolean Lombiq.Unum.Unum::IsPositive().0
                case \Hast::InternalInvocationProxy().Unum::get_SignBitMask().Unum::IsPositive().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::IsPositive().0.Unum::get_SignBitMask()._Started.0\) then 
                            \Unum::IsPositive().0.Unum::get_SignBitMask()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::get_SignBitMask().Unum::IsPositive().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::get_SignBitMask().Unum::IsPositive().0.runningIndex.0\ := 0;
                            \Unum::get_SignBitMask().0._Started\ <= true;
                            \Unum::get_SignBitMask().0.this.parameter.In\ <= \Unum::IsPositive().0.Unum::get_SignBitMask().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::get_SignBitMask().Unum::IsPositive().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::get_SignBitMask().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::get_SignBitMask().Unum::IsPositive().0.runningState.0\ := AfterFinished;
                                    \Unum::IsPositive().0.Unum::get_SignBitMask()._Finished.0\ <= true;
                                    \Unum::get_SignBitMask().0._Started\ <= false;
                                    \Unum::IsPositive().0.Unum::get_SignBitMask().return.0\ <= \Unum::get_SignBitMask().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::IsPositive().0.Unum::get_SignBitMask()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::get_SignBitMask().Unum::IsPositive().0.runningState.0\ := WaitingForStarted;
                            \Unum::IsPositive().0.Unum::get_SignBitMask()._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_SignBitMask() end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit() start
    \Hast::InternalInvocationProxy().Unum::FractionWithHiddenBit()\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Unum::FractionWithHiddenBit().Unum::FractionToUintArray().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::FractionWithHiddenBit().Unum::FractionToUintArray().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Unum::FractionWithHiddenBit().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::FractionWithHiddenBit().Unum::AddExactUnums(Unum,Unum).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().Unum::FractionWithHiddenBit().Unum::FractionToUintArray().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::FractionWithHiddenBit().Unum::FractionToUintArray().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Unum::FractionWithHiddenBit().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::FractionWithHiddenBit().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                \Unum::FractionToUintArray().0.Unum::FractionWithHiddenBit()._Finished.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.UInt32[] Lombiq.Unum.Unum::FractionToUintArray().0
                case \Hast::InternalInvocationProxy().Unum::FractionWithHiddenBit().Unum::FractionToUintArray().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::FractionToUintArray().0.Unum::FractionWithHiddenBit()._Started.0\) then 
                            \Unum::FractionToUintArray().0.Unum::FractionWithHiddenBit()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::FractionWithHiddenBit().Unum::FractionToUintArray().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::FractionWithHiddenBit().Unum::FractionToUintArray().0.runningIndex.0\ := 0;
                            \Unum::FractionWithHiddenBit().0._Started\ <= true;
                            \Unum::FractionWithHiddenBit().0.this.parameter.In\ <= \Unum::FractionToUintArray().0.Unum::FractionWithHiddenBit().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::FractionWithHiddenBit().Unum::FractionToUintArray().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::FractionWithHiddenBit().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::FractionWithHiddenBit().Unum::FractionToUintArray().0.runningState.0\ := AfterFinished;
                                    \Unum::FractionToUintArray().0.Unum::FractionWithHiddenBit()._Finished.0\ <= true;
                                    \Unum::FractionWithHiddenBit().0._Started\ <= false;
                                    \Unum::FractionToUintArray().0.Unum::FractionWithHiddenBit().return.0\ <= \Unum::FractionWithHiddenBit().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::FractionToUintArray().0.Unum::FractionWithHiddenBit()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::FractionWithHiddenBit().Unum::FractionToUintArray().0.runningState.0\ := WaitingForStarted;
                            \Unum::FractionToUintArray().0.Unum::FractionWithHiddenBit()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0
                case \Hast::InternalInvocationProxy().Unum::FractionWithHiddenBit().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Started.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::FractionWithHiddenBit().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::FractionWithHiddenBit().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                            \Unum::FractionWithHiddenBit().0._Started\ <= true;
                            \Unum::FractionWithHiddenBit().0.this.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::FractionWithHiddenBit().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::FractionWithHiddenBit().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::FractionWithHiddenBit().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := AfterFinished;
                                    \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Finished.0\ <= true;
                                    \Unum::FractionWithHiddenBit().0._Started\ <= false;
                                    \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit().return.0\ <= \Unum::FractionWithHiddenBit().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::FractionWithHiddenBit().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionWithHiddenBit()._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit() end


    -- System.Void Hast::InternalInvocationProxy().System.Int32 Lombiq.Unum.Unum::ExponentValueWithBias() start
    \Hast::InternalInvocationProxy().Unum::ExponentValueWithBias()\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Unum::ExponentValueWithBias().Unum::FractionToUintArray().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::ExponentValueWithBias().Unum::FractionToUintArray().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Unum::ExponentValueWithBias().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::ExponentValueWithBias().Unum::AddExactUnums(Unum,Unum).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().Unum::ExponentValueWithBias().Unum::FractionToUintArray().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::ExponentValueWithBias().Unum::FractionToUintArray().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Unum::ExponentValueWithBias().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::ExponentValueWithBias().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                \Unum::FractionToUintArray().0.Unum::ExponentValueWithBias()._Finished.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.UInt32[] Lombiq.Unum.Unum::FractionToUintArray().0
                case \Hast::InternalInvocationProxy().Unum::ExponentValueWithBias().Unum::FractionToUintArray().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::FractionToUintArray().0.Unum::ExponentValueWithBias()._Started.0\) then 
                            \Unum::FractionToUintArray().0.Unum::ExponentValueWithBias()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::ExponentValueWithBias().Unum::FractionToUintArray().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::ExponentValueWithBias().Unum::FractionToUintArray().0.runningIndex.0\ := 0;
                            \Unum::ExponentValueWithBias().0._Started\ <= true;
                            \Unum::ExponentValueWithBias().0.this.parameter.In\ <= \Unum::FractionToUintArray().0.Unum::ExponentValueWithBias().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::ExponentValueWithBias().Unum::FractionToUintArray().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::ExponentValueWithBias().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::ExponentValueWithBias().Unum::FractionToUintArray().0.runningState.0\ := AfterFinished;
                                    \Unum::FractionToUintArray().0.Unum::ExponentValueWithBias()._Finished.0\ <= true;
                                    \Unum::ExponentValueWithBias().0._Started\ <= false;
                                    \Unum::FractionToUintArray().0.Unum::ExponentValueWithBias().return.0\ <= \Unum::ExponentValueWithBias().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::FractionToUintArray().0.Unum::ExponentValueWithBias()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::ExponentValueWithBias().Unum::FractionToUintArray().0.runningState.0\ := WaitingForStarted;
                            \Unum::FractionToUintArray().0.Unum::ExponentValueWithBias()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0
                case \Hast::InternalInvocationProxy().Unum::ExponentValueWithBias().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Started.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::ExponentValueWithBias().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::ExponentValueWithBias().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                            \Unum::ExponentValueWithBias().0._Started\ <= true;
                            \Unum::ExponentValueWithBias().0.this.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::ExponentValueWithBias().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::ExponentValueWithBias().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::ExponentValueWithBias().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := AfterFinished;
                                    \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Finished.0\ <= true;
                                    \Unum::ExponentValueWithBias().0._Started\ <= false;
                                    \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias().return.0\ <= \Unum::ExponentValueWithBias().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::ExponentValueWithBias().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueWithBias()._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.Int32 Lombiq.Unum.Unum::ExponentValueWithBias() end


    -- System.Void Hast::InternalInvocationProxy().System.UInt16 Lombiq.Unum.Unum::FractionSize() start
    \Hast::InternalInvocationProxy().Unum::FractionSize()\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionToUintArray().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionToUintArray().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionMask().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionMask().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::ExponentMask().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::ExponentMask().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::Exponent().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::Exponent().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionWithHiddenBit().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionWithHiddenBit().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::AddExactUnums(Unum,Unum).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionToUintArray().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionToUintArray().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionMask().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionMask().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::ExponentMask().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::ExponentMask().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::Exponent().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::Exponent().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionWithHiddenBit().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionWithHiddenBit().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                \Unum::FractionToUintArray().0.Unum::FractionSize()._Finished.0\ <= false;
                \Unum::FractionMask().0.Unum::FractionSize()._Finished.0\ <= false;
                \Unum::ExponentMask().0.Unum::FractionSize()._Finished.0\ <= false;
                \Unum::Exponent().0.Unum::FractionSize()._Finished.0\ <= false;
                \Unum::FractionWithHiddenBit().0.Unum::FractionSize()._Finished.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.UInt32[] Lombiq.Unum.Unum::FractionToUintArray().0
                case \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionToUintArray().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::FractionToUintArray().0.Unum::FractionSize()._Started.0\) then 
                            \Unum::FractionToUintArray().0.Unum::FractionSize()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionToUintArray().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionToUintArray().0.runningIndex.0\ := 0;
                            \Unum::FractionSize().0._Started\ <= true;
                            \Unum::FractionSize().0.this.parameter.In\ <= \Unum::FractionToUintArray().0.Unum::FractionSize().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionToUintArray().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::FractionSize().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionToUintArray().0.runningState.0\ := AfterFinished;
                                    \Unum::FractionToUintArray().0.Unum::FractionSize()._Finished.0\ <= true;
                                    \Unum::FractionSize().0._Started\ <= false;
                                    \Unum::FractionToUintArray().0.Unum::FractionSize().return.0\ <= \Unum::FractionSize().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::FractionToUintArray().0.Unum::FractionSize()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionToUintArray().0.runningState.0\ := WaitingForStarted;
                            \Unum::FractionToUintArray().0.Unum::FractionSize()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionMask().0
                case \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionMask().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::FractionMask().0.Unum::FractionSize()._Started.0\) then 
                            \Unum::FractionMask().0.Unum::FractionSize()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionMask().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionMask().0.runningIndex.0\ := 0;
                            \Unum::FractionSize().0._Started\ <= true;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionMask().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::FractionSize().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionMask().0.runningState.0\ := AfterFinished;
                                    \Unum::FractionMask().0.Unum::FractionSize()._Finished.0\ <= true;
                                    \Unum::FractionSize().0._Started\ <= false;
                                    \Unum::FractionMask().0.Unum::FractionSize().return.0\ <= \Unum::FractionSize().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::FractionMask().0.Unum::FractionSize()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionMask().0.runningState.0\ := WaitingForStarted;
                            \Unum::FractionMask().0.Unum::FractionSize()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentMask().0
                case \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::ExponentMask().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::ExponentMask().0.Unum::FractionSize()._Started.0\) then 
                            \Unum::ExponentMask().0.Unum::FractionSize()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::ExponentMask().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::ExponentMask().0.runningIndex.0\ := 0;
                            \Unum::FractionSize().0._Started\ <= true;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::ExponentMask().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::FractionSize().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::ExponentMask().0.runningState.0\ := AfterFinished;
                                    \Unum::ExponentMask().0.Unum::FractionSize()._Finished.0\ <= true;
                                    \Unum::FractionSize().0._Started\ <= false;
                                    \Unum::ExponentMask().0.Unum::FractionSize().return.0\ <= \Unum::FractionSize().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::ExponentMask().0.Unum::FractionSize()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::ExponentMask().0.runningState.0\ := WaitingForStarted;
                            \Unum::ExponentMask().0.Unum::FractionSize()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::Exponent().0
                case \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::Exponent().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::Exponent().0.Unum::FractionSize()._Started.0\) then 
                            \Unum::Exponent().0.Unum::FractionSize()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::Exponent().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::Exponent().0.runningIndex.0\ := 0;
                            \Unum::FractionSize().0._Started\ <= true;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::Exponent().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::FractionSize().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::Exponent().0.runningState.0\ := AfterFinished;
                                    \Unum::Exponent().0.Unum::FractionSize()._Finished.0\ <= true;
                                    \Unum::FractionSize().0._Started\ <= false;
                                    \Unum::Exponent().0.Unum::FractionSize().return.0\ <= \Unum::FractionSize().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::Exponent().0.Unum::FractionSize()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::Exponent().0.runningState.0\ := WaitingForStarted;
                            \Unum::Exponent().0.Unum::FractionSize()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit().0
                case \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionWithHiddenBit().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::FractionWithHiddenBit().0.Unum::FractionSize()._Started.0\) then 
                            \Unum::FractionWithHiddenBit().0.Unum::FractionSize()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionWithHiddenBit().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionWithHiddenBit().0.runningIndex.0\ := 0;
                            \Unum::FractionSize().0._Started\ <= true;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionWithHiddenBit().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::FractionSize().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionWithHiddenBit().0.runningState.0\ := AfterFinished;
                                    \Unum::FractionWithHiddenBit().0.Unum::FractionSize()._Finished.0\ <= true;
                                    \Unum::FractionSize().0._Started\ <= false;
                                    \Unum::FractionWithHiddenBit().0.Unum::FractionSize().return.0\ <= \Unum::FractionSize().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::FractionWithHiddenBit().0.Unum::FractionSize()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::FractionWithHiddenBit().0.runningState.0\ := WaitingForStarted;
                            \Unum::FractionWithHiddenBit().0.Unum::FractionSize()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0
                case \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Started.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                            \Unum::FractionSize().0._Started\ <= true;
                            \Unum::FractionSize().0.this.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::FractionSize().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := AfterFinished;
                                    \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Finished.0\ <= true;
                                    \Unum::FractionSize().0._Started\ <= false;
                                    \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize().return.0\ <= \Unum::FractionSize().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::FractionSize().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::FractionSize()._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.UInt16 Lombiq.Unum.Unum::FractionSize() end


    -- System.Void Hast::InternalInvocationProxy().System.Boolean Lombiq.Unum.Unum::IsPositive() start
    \Hast::InternalInvocationProxy().Unum::IsPositive()\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Unum::IsPositive().Unum::FractionToUintArray().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::IsPositive().Unum::FractionToUintArray().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Unum::IsPositive().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::IsPositive().Unum::AddExactUnums(Unum,Unum).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().Unum::IsPositive().Unum::FractionToUintArray().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::IsPositive().Unum::FractionToUintArray().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Unum::IsPositive().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::IsPositive().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                \Unum::FractionToUintArray().0.Unum::IsPositive()._Finished.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.UInt32[] Lombiq.Unum.Unum::FractionToUintArray().0
                case \Hast::InternalInvocationProxy().Unum::IsPositive().Unum::FractionToUintArray().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::FractionToUintArray().0.Unum::IsPositive()._Started.0\) then 
                            \Unum::FractionToUintArray().0.Unum::IsPositive()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::IsPositive().Unum::FractionToUintArray().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::IsPositive().Unum::FractionToUintArray().0.runningIndex.0\ := 0;
                            \Unum::IsPositive().0._Started\ <= true;
                            \Unum::IsPositive().0.this.parameter.In\ <= \Unum::FractionToUintArray().0.Unum::IsPositive().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::IsPositive().Unum::FractionToUintArray().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::IsPositive().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::IsPositive().Unum::FractionToUintArray().0.runningState.0\ := AfterFinished;
                                    \Unum::FractionToUintArray().0.Unum::IsPositive()._Finished.0\ <= true;
                                    \Unum::IsPositive().0._Started\ <= false;
                                    \Unum::FractionToUintArray().0.Unum::IsPositive().return.0\ <= \Unum::IsPositive().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::FractionToUintArray().0.Unum::IsPositive()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::IsPositive().Unum::FractionToUintArray().0.runningState.0\ := WaitingForStarted;
                            \Unum::FractionToUintArray().0.Unum::IsPositive()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0
                case \Hast::InternalInvocationProxy().Unum::IsPositive().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::IsPositive().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::IsPositive().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                            \Unum::IsPositive().0._Started\ <= true;
                            \Unum::IsPositive().0.this.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::IsPositive().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::IsPositive().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::IsPositive().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := AfterFinished;
                                    \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Finished.0\ <= true;
                                    \Unum::IsPositive().0._Started\ <= false;
                                    \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive().return.0\ <= \Unum::IsPositive().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::IsPositive().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositive()._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.Boolean Lombiq.Unum.Unum::IsPositive() end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseAnd(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask) start
    \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::IsExact().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::IsExact().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::IsPositive().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::IsPositive().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::ExponentSize().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::ExponentSize().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::FractionSize().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::FractionSize().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::Exponent().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::Exponent().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::Fraction().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::Fraction().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::IsExact().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::IsExact().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::IsPositive().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::IsPositive().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::ExponentSize().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::ExponentSize().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::FractionSize().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::FractionSize().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::Exponent().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::Exponent().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::Fraction().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::Fraction().0.runningState.0\ := WaitingForStarted;
                \Unum::IsExact().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= false;
                \Unum::IsPositive().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= false;
                \Unum::ExponentSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= false;
                \Unum::FractionSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= false;
                \Unum::Exponent().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= false;
                \Unum::Fraction().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.Boolean Lombiq.Unum.Unum::IsExact().0
                case \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::IsExact().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::IsExact().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\) then 
                            \Unum::IsExact().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::IsExact().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::IsExact().0.runningIndex.0\ := 0;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0._Started\ <= true;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.left.parameter.In\ <= \Unum::IsExact().0.BitMask::op_BitwiseAnd(BitMask,BitMask).left.parameter.Out.0\;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.right.parameter.In\ <= \Unum::IsExact().0.BitMask::op_BitwiseAnd(BitMask,BitMask).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::IsExact().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_BitwiseAnd(BitMask,BitMask).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::IsExact().0.runningState.0\ := AfterFinished;
                                    \Unum::IsExact().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= true;
                                    \BitMask::op_BitwiseAnd(BitMask,BitMask).0._Started\ <= false;
                                    \Unum::IsExact().0.BitMask::op_BitwiseAnd(BitMask,BitMask).return.0\ <= \BitMask::op_BitwiseAnd(BitMask,BitMask).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::IsExact().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::IsExact().0.runningState.0\ := WaitingForStarted;
                            \Unum::IsExact().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Boolean Lombiq.Unum.Unum::IsPositive().0
                case \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::IsPositive().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::IsPositive().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\) then 
                            \Unum::IsPositive().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::IsPositive().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::IsPositive().0.runningIndex.0\ := 0;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0._Started\ <= true;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.left.parameter.In\ <= \Unum::IsPositive().0.BitMask::op_BitwiseAnd(BitMask,BitMask).left.parameter.Out.0\;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.right.parameter.In\ <= \Unum::IsPositive().0.BitMask::op_BitwiseAnd(BitMask,BitMask).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::IsPositive().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_BitwiseAnd(BitMask,BitMask).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::IsPositive().0.runningState.0\ := AfterFinished;
                                    \Unum::IsPositive().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= true;
                                    \BitMask::op_BitwiseAnd(BitMask,BitMask).0._Started\ <= false;
                                    \Unum::IsPositive().0.BitMask::op_BitwiseAnd(BitMask,BitMask).return.0\ <= \BitMask::op_BitwiseAnd(BitMask,BitMask).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::IsPositive().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::IsPositive().0.runningState.0\ := WaitingForStarted;
                            \Unum::IsPositive().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Byte Lombiq.Unum.Unum::ExponentSize().0
                case \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::ExponentSize().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::ExponentSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\) then 
                            \Unum::ExponentSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::ExponentSize().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::ExponentSize().0.runningIndex.0\ := 0;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0._Started\ <= true;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.left.parameter.In\ <= \Unum::ExponentSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask).left.parameter.Out.0\;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.right.parameter.In\ <= \Unum::ExponentSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::ExponentSize().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_BitwiseAnd(BitMask,BitMask).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::ExponentSize().0.runningState.0\ := AfterFinished;
                                    \Unum::ExponentSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= true;
                                    \BitMask::op_BitwiseAnd(BitMask,BitMask).0._Started\ <= false;
                                    \Unum::ExponentSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask).return.0\ <= \BitMask::op_BitwiseAnd(BitMask,BitMask).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::ExponentSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::ExponentSize().0.runningState.0\ := WaitingForStarted;
                            \Unum::ExponentSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.UInt16 Lombiq.Unum.Unum::FractionSize().0
                case \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::FractionSize().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::FractionSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\) then 
                            \Unum::FractionSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::FractionSize().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::FractionSize().0.runningIndex.0\ := 0;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0._Started\ <= true;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.left.parameter.In\ <= \Unum::FractionSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask).left.parameter.Out.0\;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.right.parameter.In\ <= \Unum::FractionSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::FractionSize().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_BitwiseAnd(BitMask,BitMask).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::FractionSize().0.runningState.0\ := AfterFinished;
                                    \Unum::FractionSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= true;
                                    \BitMask::op_BitwiseAnd(BitMask,BitMask).0._Started\ <= false;
                                    \Unum::FractionSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask).return.0\ <= \BitMask::op_BitwiseAnd(BitMask,BitMask).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::FractionSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::FractionSize().0.runningState.0\ := WaitingForStarted;
                            \Unum::FractionSize().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::Exponent().0
                case \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::Exponent().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::Exponent().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\) then 
                            \Unum::Exponent().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::Exponent().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::Exponent().0.runningIndex.0\ := 0;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0._Started\ <= true;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.left.parameter.In\ <= \Unum::Exponent().0.BitMask::op_BitwiseAnd(BitMask,BitMask).left.parameter.Out.0\;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.right.parameter.In\ <= \Unum::Exponent().0.BitMask::op_BitwiseAnd(BitMask,BitMask).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::Exponent().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_BitwiseAnd(BitMask,BitMask).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::Exponent().0.runningState.0\ := AfterFinished;
                                    \Unum::Exponent().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= true;
                                    \BitMask::op_BitwiseAnd(BitMask,BitMask).0._Started\ <= false;
                                    \Unum::Exponent().0.BitMask::op_BitwiseAnd(BitMask,BitMask).return.0\ <= \BitMask::op_BitwiseAnd(BitMask,BitMask).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::Exponent().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::Exponent().0.runningState.0\ := WaitingForStarted;
                            \Unum::Exponent().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::Fraction().0
                case \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::Fraction().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::Fraction().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\) then 
                            \Unum::Fraction().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::Fraction().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::Fraction().0.runningIndex.0\ := 0;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0._Started\ <= true;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.left.parameter.In\ <= \Unum::Fraction().0.BitMask::op_BitwiseAnd(BitMask,BitMask).left.parameter.Out.0\;
                            \BitMask::op_BitwiseAnd(BitMask,BitMask).0.right.parameter.In\ <= \Unum::Fraction().0.BitMask::op_BitwiseAnd(BitMask,BitMask).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::Fraction().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_BitwiseAnd(BitMask,BitMask).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::Fraction().0.runningState.0\ := AfterFinished;
                                    \Unum::Fraction().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= true;
                                    \BitMask::op_BitwiseAnd(BitMask,BitMask).0._Started\ <= false;
                                    \Unum::Fraction().0.BitMask::op_BitwiseAnd(BitMask,BitMask).return.0\ <= \BitMask::op_BitwiseAnd(BitMask,BitMask).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::Fraction().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_BitwiseAnd(BitMask,BitMask).Unum::Fraction().0.runningState.0\ := WaitingForStarted;
                            \Unum::Fraction().0.BitMask::op_BitwiseAnd(BitMask,BitMask)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseAnd(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask) end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_ExponentSizeMask() start
    -- Signal connections for System.Byte Lombiq.Unum.Unum::ExponentSize().0 (#0):
    \Unum::get_ExponentSizeMask().0._Started\ <= \Unum::ExponentSize().0.Unum::get_ExponentSizeMask()._Started.0\;
    \Unum::get_ExponentSizeMask().0.this.parameter.In\ <= \Unum::ExponentSize().0.Unum::get_ExponentSizeMask().this.parameter.Out.0\;
    \Unum::ExponentSize().0.Unum::get_ExponentSizeMask()._Finished.0\ <= \Unum::get_ExponentSizeMask().0._Finished\;
    \Unum::ExponentSize().0.Unum::get_ExponentSizeMask().return.0\ <= \Unum::get_ExponentSizeMask().0.return\;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_ExponentSizeMask() end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_FractionSizeMask() start
    -- Signal connections for System.UInt16 Lombiq.Unum.Unum::FractionSize().0 (#0):
    \Unum::get_FractionSizeMask().0._Started\ <= \Unum::FractionSize().0.Unum::get_FractionSizeMask()._Started.0\;
    \Unum::get_FractionSizeMask().0.this.parameter.In\ <= \Unum::FractionSize().0.Unum::get_FractionSizeMask().this.parameter.Out.0\;
    \Unum::FractionSize().0.Unum::get_FractionSizeMask()._Finished.0\ <= \Unum::get_FractionSizeMask().0._Finished\;
    \Unum::FractionSize().0.Unum::get_FractionSizeMask().return.0\ <= \Unum::get_FractionSizeMask().0.return\;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_FractionSizeMask() end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,System.UInt32) start
    \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::FractionMask().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::FractionMask().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::ExponentMask().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::ExponentMask().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::FractionMask().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::FractionMask().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::ExponentMask().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::ExponentMask().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := WaitingForStarted;
                \Unum::FractionMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\ <= false;
                \Unum::ExponentMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\ <= false;
                \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\ <= false;
                \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionMask().0
                case \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::FractionMask().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::FractionMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\) then 
                            \Unum::FractionMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::FractionMask().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::FractionMask().0.runningIndex.0\ := 0;
                            \BitMask::op_Subtraction(BitMask,UInt32).0._Started\ <= true;
                            \BitMask::op_Subtraction(BitMask,UInt32).0.left.parameter.In\ <= \Unum::FractionMask().0.BitMask::op_Subtraction(BitMask,UInt32).left.parameter.Out.0\;
                            \BitMask::op_Subtraction(BitMask,UInt32).0.right.parameter.In\ <= \Unum::FractionMask().0.BitMask::op_Subtraction(BitMask,UInt32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::FractionMask().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Subtraction(BitMask,UInt32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::FractionMask().0.runningState.0\ := AfterFinished;
                                    \Unum::FractionMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\ <= true;
                                    \BitMask::op_Subtraction(BitMask,UInt32).0._Started\ <= false;
                                    \Unum::FractionMask().0.BitMask::op_Subtraction(BitMask,UInt32).return.0\ <= \BitMask::op_Subtraction(BitMask,UInt32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::FractionMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::FractionMask().0.runningState.0\ := WaitingForStarted;
                            \Unum::FractionMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentMask().0
                case \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::ExponentMask().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::ExponentMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\) then 
                            \Unum::ExponentMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::ExponentMask().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::ExponentMask().0.runningIndex.0\ := 0;
                            \BitMask::op_Subtraction(BitMask,UInt32).0._Started\ <= true;
                            \BitMask::op_Subtraction(BitMask,UInt32).0.left.parameter.In\ <= \Unum::ExponentMask().0.BitMask::op_Subtraction(BitMask,UInt32).left.parameter.Out.0\;
                            \BitMask::op_Subtraction(BitMask,UInt32).0.right.parameter.In\ <= \Unum::ExponentMask().0.BitMask::op_Subtraction(BitMask,UInt32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::ExponentMask().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Subtraction(BitMask,UInt32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::ExponentMask().0.runningState.0\ := AfterFinished;
                                    \Unum::ExponentMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\ <= true;
                                    \BitMask::op_Subtraction(BitMask,UInt32).0._Started\ <= false;
                                    \Unum::ExponentMask().0.BitMask::op_Subtraction(BitMask,UInt32).return.0\ <= \BitMask::op_Subtraction(BitMask,UInt32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::ExponentMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::ExponentMask().0.runningState.0\ := WaitingForStarted;
                            \Unum::ExponentMask().0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentValueToExponentBits(System.Int32,System.Byte).0
                case \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\) then 
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningIndex.0\ := 0;
                            \BitMask::op_Subtraction(BitMask,UInt32).0._Started\ <= true;
                            \BitMask::op_Subtraction(BitMask,UInt32).0.left.parameter.In\ <= \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).left.parameter.Out.0\;
                            \BitMask::op_Subtraction(BitMask,UInt32).0.right.parameter.In\ <= \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Subtraction(BitMask,UInt32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningState.0\ := AfterFinished;
                                    \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\ <= true;
                                    \BitMask::op_Subtraction(BitMask,UInt32).0._Started\ <= false;
                                    \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).return.0\ <= \BitMask::op_Subtraction(BitMask,UInt32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).Unum::ExponentValueToExponentBits(Int32,Byte).0.runningState.0\ := WaitingForStarted;
                            \Unum::ExponentValueToExponentBits(Int32,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Void Lombiq.Unum.UnumEnvironment::.ctor(System.Byte,System.Byte).0
                case \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\ := 0;
                            \BitMask::op_Subtraction(BitMask,UInt32).0._Started\ <= true;
                            \BitMask::op_Subtraction(BitMask,UInt32).0.left.parameter.In\ <= \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).left.parameter.Out.0\;
                            \BitMask::op_Subtraction(BitMask,UInt32).0.right.parameter.In\ <= \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::op_Subtraction(BitMask,UInt32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := AfterFinished;
                                    \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\ <= true;
                                    \BitMask::op_Subtraction(BitMask,UInt32).0._Started\ <= false;
                                    \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32).return.0\ <= \BitMask::op_Subtraction(BitMask,UInt32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::op_Subtraction(BitMask,UInt32).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := WaitingForStarted;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_Subtraction(BitMask,UInt32)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_Subtraction(Lombiq.Unum.BitMask,System.UInt32) end


    -- System.Void Hast::InternalInvocationProxy().System.Byte Lombiq.Unum.Unum::ExponentSize() start
    \Hast::InternalInvocationProxy().Unum::ExponentSize()\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Unum::ExponentSize().Unum::ExponentMask().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::ExponentSize().Unum::ExponentMask().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Unum::ExponentSize().Unum::Bias().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::ExponentSize().Unum::Bias().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().Unum::ExponentSize().Unum::ExponentMask().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::ExponentSize().Unum::ExponentMask().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Unum::ExponentSize().Unum::Bias().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::ExponentSize().Unum::Bias().0.runningState.0\ := WaitingForStarted;
                \Unum::ExponentMask().0.Unum::ExponentSize()._Finished.0\ <= false;
                \Unum::Bias().0.Unum::ExponentSize()._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentMask().0
                case \Hast::InternalInvocationProxy().Unum::ExponentSize().Unum::ExponentMask().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::ExponentMask().0.Unum::ExponentSize()._Started.0\) then 
                            \Unum::ExponentMask().0.Unum::ExponentSize()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::ExponentSize().Unum::ExponentMask().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::ExponentSize().Unum::ExponentMask().0.runningIndex.0\ := 0;
                            \Unum::ExponentSize().0._Started\ <= true;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::ExponentSize().Unum::ExponentMask().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::ExponentSize().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::ExponentSize().Unum::ExponentMask().0.runningState.0\ := AfterFinished;
                                    \Unum::ExponentMask().0.Unum::ExponentSize()._Finished.0\ <= true;
                                    \Unum::ExponentSize().0._Started\ <= false;
                                    \Unum::ExponentMask().0.Unum::ExponentSize().return.0\ <= \Unum::ExponentSize().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::ExponentMask().0.Unum::ExponentSize()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::ExponentSize().Unum::ExponentMask().0.runningState.0\ := WaitingForStarted;
                            \Unum::ExponentMask().0.Unum::ExponentSize()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Int32 Lombiq.Unum.Unum::Bias().0
                case \Hast::InternalInvocationProxy().Unum::ExponentSize().Unum::Bias().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::Bias().0.Unum::ExponentSize()._Started.0\) then 
                            \Unum::Bias().0.Unum::ExponentSize()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::ExponentSize().Unum::Bias().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::ExponentSize().Unum::Bias().0.runningIndex.0\ := 0;
                            \Unum::ExponentSize().0._Started\ <= true;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::ExponentSize().Unum::Bias().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::ExponentSize().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::ExponentSize().Unum::Bias().0.runningState.0\ := AfterFinished;
                                    \Unum::Bias().0.Unum::ExponentSize()._Finished.0\ <= true;
                                    \Unum::ExponentSize().0._Started\ <= false;
                                    \Unum::Bias().0.Unum::ExponentSize().return.0\ <= \Unum::ExponentSize().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::Bias().0.Unum::ExponentSize()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::ExponentSize().Unum::Bias().0.runningState.0\ := WaitingForStarted;
                            \Unum::Bias().0.Unum::ExponentSize()._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.Byte Lombiq.Unum.Unum::ExponentSize() end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentMask() start
    -- Signal connections for Lombiq.Unum.BitMask Lombiq.Unum.Unum::Exponent().0 (#0):
    \Unum::ExponentMask().0._Started\ <= \Unum::Exponent().0.Unum::ExponentMask()._Started.0\;
    \Unum::Exponent().0.Unum::ExponentMask()._Finished.0\ <= \Unum::ExponentMask().0._Finished\;
    \Unum::Exponent().0.Unum::ExponentMask().return.0\ <= \Unum::ExponentMask().0.return\;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentMask() end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionMask() start
    -- Signal connections for Lombiq.Unum.BitMask Lombiq.Unum.Unum::Fraction().0 (#0):
    \Unum::FractionMask().0._Started\ <= \Unum::Fraction().0.Unum::FractionMask()._Started.0\;
    \Unum::Fraction().0.Unum::FractionMask()._Finished.0\ <= \Unum::FractionMask().0._Finished\;
    \Unum::Fraction().0.Unum::FractionMask().return.0\ <= \Unum::FractionMask().0.return\;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionMask() end


    -- System.Void Hast::InternalInvocationProxy().System.Boolean Lombiq.Unum.Unum::HiddenBitIsOne() start
    \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne()\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::FractionWithHiddenBit().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::FractionWithHiddenBit().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::ExponentValueWithBias().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::ExponentValueWithBias().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::AddExactUnums(Unum,Unum).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::FractionWithHiddenBit().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::FractionWithHiddenBit().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::ExponentValueWithBias().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::ExponentValueWithBias().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                \Unum::FractionWithHiddenBit().0.Unum::HiddenBitIsOne()._Finished.0\ <= false;
                \Unum::ExponentValueWithBias().0.Unum::HiddenBitIsOne()._Finished.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne()._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit().0
                case \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::FractionWithHiddenBit().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::FractionWithHiddenBit().0.Unum::HiddenBitIsOne()._Started.0\) then 
                            \Unum::FractionWithHiddenBit().0.Unum::HiddenBitIsOne()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::FractionWithHiddenBit().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::FractionWithHiddenBit().0.runningIndex.0\ := 0;
                            \Unum::HiddenBitIsOne().0._Started\ <= true;
                            \Unum::HiddenBitIsOne().0.this.parameter.In\ <= \Unum::FractionWithHiddenBit().0.Unum::HiddenBitIsOne().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::FractionWithHiddenBit().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::HiddenBitIsOne().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::FractionWithHiddenBit().0.runningState.0\ := AfterFinished;
                                    \Unum::FractionWithHiddenBit().0.Unum::HiddenBitIsOne()._Finished.0\ <= true;
                                    \Unum::HiddenBitIsOne().0._Started\ <= false;
                                    \Unum::FractionWithHiddenBit().0.Unum::HiddenBitIsOne().return.0\ <= \Unum::HiddenBitIsOne().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::FractionWithHiddenBit().0.Unum::HiddenBitIsOne()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::FractionWithHiddenBit().0.runningState.0\ := WaitingForStarted;
                            \Unum::FractionWithHiddenBit().0.Unum::HiddenBitIsOne()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Int32 Lombiq.Unum.Unum::ExponentValueWithBias().0
                case \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::ExponentValueWithBias().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::ExponentValueWithBias().0.Unum::HiddenBitIsOne()._Started.0\) then 
                            \Unum::ExponentValueWithBias().0.Unum::HiddenBitIsOne()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::ExponentValueWithBias().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::ExponentValueWithBias().0.runningIndex.0\ := 0;
                            \Unum::HiddenBitIsOne().0._Started\ <= true;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::ExponentValueWithBias().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::HiddenBitIsOne().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::ExponentValueWithBias().0.runningState.0\ := AfterFinished;
                                    \Unum::ExponentValueWithBias().0.Unum::HiddenBitIsOne()._Finished.0\ <= true;
                                    \Unum::HiddenBitIsOne().0._Started\ <= false;
                                    \Unum::ExponentValueWithBias().0.Unum::HiddenBitIsOne().return.0\ <= \Unum::HiddenBitIsOne().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::ExponentValueWithBias().0.Unum::HiddenBitIsOne()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::ExponentValueWithBias().0.runningState.0\ := WaitingForStarted;
                            \Unum::ExponentValueWithBias().0.Unum::HiddenBitIsOne()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0
                case \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne()._Started.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                            \Unum::HiddenBitIsOne().0._Started\ <= true;
                            \Unum::HiddenBitIsOne().0.this.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::HiddenBitIsOne().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := AfterFinished;
                                    \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne()._Finished.0\ <= true;
                                    \Unum::HiddenBitIsOne().0._Started\ <= false;
                                    \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne().return.0\ <= \Unum::HiddenBitIsOne().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::HiddenBitIsOne().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::HiddenBitIsOne()._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.Boolean Lombiq.Unum.Unum::HiddenBitIsOne() end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::Fraction() start
    \Hast::InternalInvocationProxy().Unum::Fraction()\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Unum::Fraction().Unum::FractionWithHiddenBit().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::Fraction().Unum::FractionWithHiddenBit().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Unum::Fraction().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::Fraction().Unum::AddExactUnums(Unum,Unum).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().Unum::Fraction().Unum::FractionWithHiddenBit().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::Fraction().Unum::FractionWithHiddenBit().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Unum::Fraction().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::Fraction().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                \Unum::FractionWithHiddenBit().0.Unum::Fraction()._Finished.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction()._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit().0
                case \Hast::InternalInvocationProxy().Unum::Fraction().Unum::FractionWithHiddenBit().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::FractionWithHiddenBit().0.Unum::Fraction()._Started.0\) then 
                            \Unum::FractionWithHiddenBit().0.Unum::Fraction()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::Fraction().Unum::FractionWithHiddenBit().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::Fraction().Unum::FractionWithHiddenBit().0.runningIndex.0\ := 0;
                            \Unum::Fraction().0._Started\ <= true;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::Fraction().Unum::FractionWithHiddenBit().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::Fraction().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::Fraction().Unum::FractionWithHiddenBit().0.runningState.0\ := AfterFinished;
                                    \Unum::FractionWithHiddenBit().0.Unum::Fraction()._Finished.0\ <= true;
                                    \Unum::Fraction().0._Started\ <= false;
                                    \Unum::FractionWithHiddenBit().0.Unum::Fraction().return.0\ <= \Unum::Fraction().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::FractionWithHiddenBit().0.Unum::Fraction()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::Fraction().Unum::FractionWithHiddenBit().0.runningState.0\ := WaitingForStarted;
                            \Unum::FractionWithHiddenBit().0.Unum::Fraction()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0
                case \Hast::InternalInvocationProxy().Unum::Fraction().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction()._Started.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::Fraction().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::Fraction().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                            \Unum::Fraction().0._Started\ <= true;
                            \Unum::Fraction().0.this.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::Fraction().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::Fraction().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::Fraction().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := AfterFinished;
                                    \Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction()._Finished.0\ <= true;
                                    \Unum::Fraction().0._Started\ <= false;
                                    \Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction().return.0\ <= \Unum::Fraction().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::Fraction().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::Fraction()._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::Fraction() end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetOne(System.UInt16) start
    \Hast::InternalInvocationProxy().BitMask::SetOne(UInt16)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().BitMask::SetOne(UInt16).Unum::FractionWithHiddenBit().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::SetOne(UInt16).Unum::FractionWithHiddenBit().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().BitMask::SetOne(UInt16).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().BitMask::SetOne(UInt16).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().BitMask::SetOne(UInt16).Unum::FractionWithHiddenBit().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::SetOne(UInt16).Unum::FractionWithHiddenBit().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().BitMask::SetOne(UInt16).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().BitMask::SetOne(UInt16).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := WaitingForStarted;
                \Unum::FractionWithHiddenBit().0.BitMask::SetOne(UInt16)._Finished.0\ <= false;
                \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.BitMask Lombiq.Unum.Unum::FractionWithHiddenBit().0
                case \Hast::InternalInvocationProxy().BitMask::SetOne(UInt16).Unum::FractionWithHiddenBit().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::FractionWithHiddenBit().0.BitMask::SetOne(UInt16)._Started.0\) then 
                            \Unum::FractionWithHiddenBit().0.BitMask::SetOne(UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::SetOne(UInt16).Unum::FractionWithHiddenBit().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::SetOne(UInt16).Unum::FractionWithHiddenBit().0.runningIndex.0\ := 0;
                            \BitMask::SetOne(UInt16).0._Started\ <= true;
                            \BitMask::SetOne(UInt16).0.this.parameter.In\ <= \Unum::FractionWithHiddenBit().0.BitMask::SetOne(UInt16).this.parameter.Out.0\;
                            \BitMask::SetOne(UInt16).0.index.parameter.In\ <= \Unum::FractionWithHiddenBit().0.BitMask::SetOne(UInt16).index.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::SetOne(UInt16).Unum::FractionWithHiddenBit().0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::SetOne(UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::SetOne(UInt16).Unum::FractionWithHiddenBit().0.runningState.0\ := AfterFinished;
                                    \Unum::FractionWithHiddenBit().0.BitMask::SetOne(UInt16)._Finished.0\ <= true;
                                    \BitMask::SetOne(UInt16).0._Started\ <= false;
                                    \Unum::FractionWithHiddenBit().0.BitMask::SetOne(UInt16).return.0\ <= \BitMask::SetOne(UInt16).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::FractionWithHiddenBit().0.BitMask::SetOne(UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::SetOne(UInt16).Unum::FractionWithHiddenBit().0.runningState.0\ := WaitingForStarted;
                            \Unum::FractionWithHiddenBit().0.BitMask::SetOne(UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Void Lombiq.Unum.UnumEnvironment::.ctor(System.Byte,System.Byte).0
                case \Hast::InternalInvocationProxy().BitMask::SetOne(UInt16).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Started.0\) then 
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().BitMask::SetOne(UInt16).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().BitMask::SetOne(UInt16).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\ := 0;
                            \BitMask::SetOne(UInt16).0._Started\ <= true;
                            \BitMask::SetOne(UInt16).0.this.parameter.In\ <= \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).this.parameter.Out.0\;
                            \BitMask::SetOne(UInt16).0.index.parameter.In\ <= \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).index.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().BitMask::SetOne(UInt16).UnumEnvironment::.ctor(Byte,Byte).0.runningIndex.0\ is 
                            when 0 => 
                                if (\BitMask::SetOne(UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().BitMask::SetOne(UInt16).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := AfterFinished;
                                    \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Finished.0\ <= true;
                                    \BitMask::SetOne(UInt16).0._Started\ <= false;
                                    \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16).return.0\ <= \BitMask::SetOne(UInt16).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().BitMask::SetOne(UInt16).UnumEnvironment::.ctor(Byte,Byte).0.runningState.0\ := WaitingForStarted;
                            \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::SetOne(UInt16)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::SetOne(System.UInt16) end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::Exponent() start
    \Hast::InternalInvocationProxy().Unum::Exponent()\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Unum::Exponent().Unum::HiddenBitIsOne().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::Exponent().Unum::HiddenBitIsOne().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Unum::Exponent().Unum::ExponentValueWithBias().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::Exponent().Unum::ExponentValueWithBias().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().Unum::Exponent().Unum::HiddenBitIsOne().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::Exponent().Unum::HiddenBitIsOne().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Unum::Exponent().Unum::ExponentValueWithBias().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::Exponent().Unum::ExponentValueWithBias().0.runningState.0\ := WaitingForStarted;
                \Unum::HiddenBitIsOne().0.Unum::Exponent()._Finished.0\ <= false;
                \Unum::ExponentValueWithBias().0.Unum::Exponent()._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.Boolean Lombiq.Unum.Unum::HiddenBitIsOne().0
                case \Hast::InternalInvocationProxy().Unum::Exponent().Unum::HiddenBitIsOne().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::HiddenBitIsOne().0.Unum::Exponent()._Started.0\) then 
                            \Unum::HiddenBitIsOne().0.Unum::Exponent()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::Exponent().Unum::HiddenBitIsOne().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::Exponent().Unum::HiddenBitIsOne().0.runningIndex.0\ := 0;
                            \Unum::Exponent().0._Started\ <= true;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::Exponent().Unum::HiddenBitIsOne().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::Exponent().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::Exponent().Unum::HiddenBitIsOne().0.runningState.0\ := AfterFinished;
                                    \Unum::HiddenBitIsOne().0.Unum::Exponent()._Finished.0\ <= true;
                                    \Unum::Exponent().0._Started\ <= false;
                                    \Unum::HiddenBitIsOne().0.Unum::Exponent().return.0\ <= \Unum::Exponent().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::HiddenBitIsOne().0.Unum::Exponent()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::Exponent().Unum::HiddenBitIsOne().0.runningState.0\ := WaitingForStarted;
                            \Unum::HiddenBitIsOne().0.Unum::Exponent()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Int32 Lombiq.Unum.Unum::ExponentValueWithBias().0
                case \Hast::InternalInvocationProxy().Unum::Exponent().Unum::ExponentValueWithBias().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::ExponentValueWithBias().0.Unum::Exponent()._Started.0\) then 
                            \Unum::ExponentValueWithBias().0.Unum::Exponent()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::Exponent().Unum::ExponentValueWithBias().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::Exponent().Unum::ExponentValueWithBias().0.runningIndex.0\ := 0;
                            \Unum::Exponent().0._Started\ <= true;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::Exponent().Unum::ExponentValueWithBias().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::Exponent().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::Exponent().Unum::ExponentValueWithBias().0.runningState.0\ := AfterFinished;
                                    \Unum::ExponentValueWithBias().0.Unum::Exponent()._Finished.0\ <= true;
                                    \Unum::Exponent().0._Started\ <= false;
                                    \Unum::ExponentValueWithBias().0.Unum::Exponent().return.0\ <= \Unum::Exponent().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::ExponentValueWithBias().0.Unum::Exponent()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::Exponent().Unum::ExponentValueWithBias().0.runningState.0\ := WaitingForStarted;
                            \Unum::ExponentValueWithBias().0.Unum::Exponent()._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::Exponent() end


    -- System.Void Hast::InternalInvocationProxy().System.Int32 Lombiq.Unum.Unum::Bias() start
    -- Signal connections for System.Int32 Lombiq.Unum.Unum::ExponentValueWithBias().0 (#0):
    \Unum::Bias().0._Started\ <= \Unum::ExponentValueWithBias().0.Unum::Bias()._Started.0\;
    \Unum::ExponentValueWithBias().0.Unum::Bias()._Finished.0\ <= \Unum::Bias().0._Finished\;
    \Unum::ExponentValueWithBias().0.Unum::Bias().return.0\ <= \Unum::Bias().0.return\;
    -- System.Void Hast::InternalInvocationProxy().System.Int32 Lombiq.Unum.Unum::Bias() end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_SignalingNotANumber() start
    -- Signal connections for System.Boolean Lombiq.Unum.Unum::IsNan().0 (#0):
    \Unum::get_SignalingNotANumber().0._Started\ <= \Unum::IsNan().0.Unum::get_SignalingNotANumber()._Started.0\;
    \Unum::get_SignalingNotANumber().0.this.parameter.In\ <= \Unum::IsNan().0.Unum::get_SignalingNotANumber().this.parameter.Out.0\;
    \Unum::IsNan().0.Unum::get_SignalingNotANumber()._Finished.0\ <= \Unum::get_SignalingNotANumber().0._Finished\;
    \Unum::IsNan().0.Unum::get_SignalingNotANumber().return.0\ <= \Unum::get_SignalingNotANumber().0.return\;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_SignalingNotANumber() end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_QuietNotANumber() start
    \Hast::InternalInvocationProxy().Unum::get_QuietNotANumber()\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Unum::get_QuietNotANumber().Unum::IsNan().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::get_QuietNotANumber().Unum::IsNan().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Unum::get_QuietNotANumber().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::get_QuietNotANumber().Unum::AddExactUnums(Unum,Unum).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().Unum::get_QuietNotANumber().Unum::IsNan().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::get_QuietNotANumber().Unum::IsNan().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Unum::get_QuietNotANumber().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::get_QuietNotANumber().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                \Unum::IsNan().0.Unum::get_QuietNotANumber()._Finished.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber()._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.Boolean Lombiq.Unum.Unum::IsNan().0
                case \Hast::InternalInvocationProxy().Unum::get_QuietNotANumber().Unum::IsNan().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::IsNan().0.Unum::get_QuietNotANumber()._Started.0\) then 
                            \Unum::IsNan().0.Unum::get_QuietNotANumber()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::get_QuietNotANumber().Unum::IsNan().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::get_QuietNotANumber().Unum::IsNan().0.runningIndex.0\ := 0;
                            \Unum::get_QuietNotANumber().0._Started\ <= true;
                            \Unum::get_QuietNotANumber().0.this.parameter.In\ <= \Unum::IsNan().0.Unum::get_QuietNotANumber().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::get_QuietNotANumber().Unum::IsNan().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::get_QuietNotANumber().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::get_QuietNotANumber().Unum::IsNan().0.runningState.0\ := AfterFinished;
                                    \Unum::IsNan().0.Unum::get_QuietNotANumber()._Finished.0\ <= true;
                                    \Unum::get_QuietNotANumber().0._Started\ <= false;
                                    \Unum::IsNan().0.Unum::get_QuietNotANumber().return.0\ <= \Unum::get_QuietNotANumber().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::IsNan().0.Unum::get_QuietNotANumber()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::get_QuietNotANumber().Unum::IsNan().0.runningState.0\ := WaitingForStarted;
                            \Unum::IsNan().0.Unum::get_QuietNotANumber()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0
                case \Hast::InternalInvocationProxy().Unum::get_QuietNotANumber().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber()._Started.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::get_QuietNotANumber().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::get_QuietNotANumber().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                            \Unum::get_QuietNotANumber().0._Started\ <= true;
                            \Unum::get_QuietNotANumber().0.this.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::get_QuietNotANumber().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::get_QuietNotANumber().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::get_QuietNotANumber().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := AfterFinished;
                                    \Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber()._Finished.0\ <= true;
                                    \Unum::get_QuietNotANumber().0._Started\ <= false;
                                    \Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber().return.0\ <= \Unum::get_QuietNotANumber().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::get_QuietNotANumber().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_QuietNotANumber()._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_QuietNotANumber() end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_PositiveInfinity() start
    \Hast::InternalInvocationProxy().Unum::get_PositiveInfinity()\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Unum::get_PositiveInfinity().Unum::IsPositiveInfinity().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::get_PositiveInfinity().Unum::IsPositiveInfinity().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Unum::get_PositiveInfinity().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::get_PositiveInfinity().Unum::AddExactUnums(Unum,Unum).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().Unum::get_PositiveInfinity().Unum::IsPositiveInfinity().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::get_PositiveInfinity().Unum::IsPositiveInfinity().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Unum::get_PositiveInfinity().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::get_PositiveInfinity().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                \Unum::IsPositiveInfinity().0.Unum::get_PositiveInfinity()._Finished.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::get_PositiveInfinity()._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.Boolean Lombiq.Unum.Unum::IsPositiveInfinity().0
                case \Hast::InternalInvocationProxy().Unum::get_PositiveInfinity().Unum::IsPositiveInfinity().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::IsPositiveInfinity().0.Unum::get_PositiveInfinity()._Started.0\) then 
                            \Unum::IsPositiveInfinity().0.Unum::get_PositiveInfinity()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::get_PositiveInfinity().Unum::IsPositiveInfinity().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::get_PositiveInfinity().Unum::IsPositiveInfinity().0.runningIndex.0\ := 0;
                            \Unum::get_PositiveInfinity().0._Started\ <= true;
                            \Unum::get_PositiveInfinity().0.this.parameter.In\ <= \Unum::IsPositiveInfinity().0.Unum::get_PositiveInfinity().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::get_PositiveInfinity().Unum::IsPositiveInfinity().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::get_PositiveInfinity().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::get_PositiveInfinity().Unum::IsPositiveInfinity().0.runningState.0\ := AfterFinished;
                                    \Unum::IsPositiveInfinity().0.Unum::get_PositiveInfinity()._Finished.0\ <= true;
                                    \Unum::get_PositiveInfinity().0._Started\ <= false;
                                    \Unum::IsPositiveInfinity().0.Unum::get_PositiveInfinity().return.0\ <= \Unum::get_PositiveInfinity().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::IsPositiveInfinity().0.Unum::get_PositiveInfinity()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::get_PositiveInfinity().Unum::IsPositiveInfinity().0.runningState.0\ := WaitingForStarted;
                            \Unum::IsPositiveInfinity().0.Unum::get_PositiveInfinity()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0
                case \Hast::InternalInvocationProxy().Unum::get_PositiveInfinity().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::get_PositiveInfinity()._Started.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_PositiveInfinity()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::get_PositiveInfinity().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::get_PositiveInfinity().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                            \Unum::get_PositiveInfinity().0._Started\ <= true;
                            \Unum::get_PositiveInfinity().0.this.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::get_PositiveInfinity().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::get_PositiveInfinity().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::get_PositiveInfinity().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::get_PositiveInfinity().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := AfterFinished;
                                    \Unum::AddExactUnums(Unum,Unum).0.Unum::get_PositiveInfinity()._Finished.0\ <= true;
                                    \Unum::get_PositiveInfinity().0._Started\ <= false;
                                    \Unum::AddExactUnums(Unum,Unum).0.Unum::get_PositiveInfinity().return.0\ <= \Unum::get_PositiveInfinity().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::get_PositiveInfinity()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::get_PositiveInfinity().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_PositiveInfinity()._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_PositiveInfinity() end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_NegativeInfinity() start
    \Hast::InternalInvocationProxy().Unum::get_NegativeInfinity()\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Unum::get_NegativeInfinity().Unum::IsNegativeInfinity().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::get_NegativeInfinity().Unum::IsNegativeInfinity().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Unum::get_NegativeInfinity().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Unum::get_NegativeInfinity().Unum::AddExactUnums(Unum,Unum).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().Unum::get_NegativeInfinity().Unum::IsNegativeInfinity().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::get_NegativeInfinity().Unum::IsNegativeInfinity().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Unum::get_NegativeInfinity().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Unum::get_NegativeInfinity().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                \Unum::IsNegativeInfinity().0.Unum::get_NegativeInfinity()._Finished.0\ <= false;
                \Unum::AddExactUnums(Unum,Unum).0.Unum::get_NegativeInfinity()._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.Boolean Lombiq.Unum.Unum::IsNegativeInfinity().0
                case \Hast::InternalInvocationProxy().Unum::get_NegativeInfinity().Unum::IsNegativeInfinity().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::IsNegativeInfinity().0.Unum::get_NegativeInfinity()._Started.0\) then 
                            \Unum::IsNegativeInfinity().0.Unum::get_NegativeInfinity()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::get_NegativeInfinity().Unum::IsNegativeInfinity().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::get_NegativeInfinity().Unum::IsNegativeInfinity().0.runningIndex.0\ := 0;
                            \Unum::get_NegativeInfinity().0._Started\ <= true;
                            \Unum::get_NegativeInfinity().0.this.parameter.In\ <= \Unum::IsNegativeInfinity().0.Unum::get_NegativeInfinity().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::get_NegativeInfinity().Unum::IsNegativeInfinity().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::get_NegativeInfinity().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::get_NegativeInfinity().Unum::IsNegativeInfinity().0.runningState.0\ := AfterFinished;
                                    \Unum::IsNegativeInfinity().0.Unum::get_NegativeInfinity()._Finished.0\ <= true;
                                    \Unum::get_NegativeInfinity().0._Started\ <= false;
                                    \Unum::IsNegativeInfinity().0.Unum::get_NegativeInfinity().return.0\ <= \Unum::get_NegativeInfinity().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::IsNegativeInfinity().0.Unum::get_NegativeInfinity()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::get_NegativeInfinity().Unum::IsNegativeInfinity().0.runningState.0\ := WaitingForStarted;
                            \Unum::IsNegativeInfinity().0.Unum::get_NegativeInfinity()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0
                case \Hast::InternalInvocationProxy().Unum::get_NegativeInfinity().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::get_NegativeInfinity()._Started.0\) then 
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_NegativeInfinity()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Unum::get_NegativeInfinity().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Unum::get_NegativeInfinity().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ := 0;
                            \Unum::get_NegativeInfinity().0._Started\ <= true;
                            \Unum::get_NegativeInfinity().0.this.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::get_NegativeInfinity().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Unum::get_NegativeInfinity().Unum::AddExactUnums(Unum,Unum).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Unum::get_NegativeInfinity().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Unum::get_NegativeInfinity().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := AfterFinished;
                                    \Unum::AddExactUnums(Unum,Unum).0.Unum::get_NegativeInfinity()._Finished.0\ <= true;
                                    \Unum::get_NegativeInfinity().0._Started\ <= false;
                                    \Unum::AddExactUnums(Unum,Unum).0.Unum::get_NegativeInfinity().return.0\ <= \Unum::get_NegativeInfinity().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Unum::AddExactUnums(Unum,Unum).0.Unum::get_NegativeInfinity()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Unum::get_NegativeInfinity().Unum::AddExactUnums(Unum,Unum).0.runningState.0\ := WaitingForStarted;
                            \Unum::AddExactUnums(Unum,Unum).0.Unum::get_NegativeInfinity()._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::get_NegativeInfinity() end


    -- System.Void Hast::InternalInvocationProxy().System.Boolean Lombiq.Unum.Unum::IsNan() start
    -- Signal connections for Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0 (#0):
    \Unum::IsNan().0._Started\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNan()._Started.0\;
    \Unum::IsNan().0.this.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNan().this.parameter.Out.0\;
    \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNan()._Finished.0\ <= \Unum::IsNan().0._Finished\;
    \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNan().return.0\ <= \Unum::IsNan().0.return\;
    -- System.Void Hast::InternalInvocationProxy().System.Boolean Lombiq.Unum.Unum::IsNan() end


    -- System.Void Hast::InternalInvocationProxy().System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,Lombiq.Unum.BitMask) start
    -- Signal connections for Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0 (#0):
    \Unum::.ctor(UnumEnvironment,BitMask).0._Started\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask)._Started.0\;
    \Unum::.ctor(UnumEnvironment,BitMask).0.this.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).this.parameter.Out.0\;
    \Unum::.ctor(UnumEnvironment,BitMask).0.environment.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).environment.parameter.Out.0\;
    \Unum::.ctor(UnumEnvironment,BitMask).0.bits.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).bits.parameter.Out.0\;
    \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask)._Finished.0\ <= \Unum::.ctor(UnumEnvironment,BitMask).0._Finished\;
    \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).this.parameter.In.0\ <= \Unum::.ctor(UnumEnvironment,BitMask).0.this.parameter.Out\;
    \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment,BitMask).environment.parameter.In.0\ <= \Unum::.ctor(UnumEnvironment,BitMask).0.environment.parameter.Out\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment,Lombiq.Unum.BitMask) end


    -- System.Void Hast::InternalInvocationProxy().System.Boolean Lombiq.Unum.Unum::IsPositiveInfinity() start
    -- Signal connections for Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0 (#0):
    \Unum::IsPositiveInfinity().0._Started\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity()._Started.0\;
    \Unum::IsPositiveInfinity().0.this.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity().this.parameter.Out.0\;
    \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity()._Finished.0\ <= \Unum::IsPositiveInfinity().0._Finished\;
    \Unum::AddExactUnums(Unum,Unum).0.Unum::IsPositiveInfinity().return.0\ <= \Unum::IsPositiveInfinity().0.return\;
    -- System.Void Hast::InternalInvocationProxy().System.Boolean Lombiq.Unum.Unum::IsPositiveInfinity() end


    -- System.Void Hast::InternalInvocationProxy().System.Boolean Lombiq.Unum.Unum::IsNegativeInfinity() start
    -- Signal connections for Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0 (#0):
    \Unum::IsNegativeInfinity().0._Started\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity()._Started.0\;
    \Unum::IsNegativeInfinity().0.this.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity().this.parameter.Out.0\;
    \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity()._Finished.0\ <= \Unum::IsNegativeInfinity().0._Finished\;
    \Unum::AddExactUnums(Unum,Unum).0.Unum::IsNegativeInfinity().return.0\ <= \Unum::IsNegativeInfinity().0.return\;
    -- System.Void Hast::InternalInvocationProxy().System.Boolean Lombiq.Unum.Unum::IsNegativeInfinity() end


    -- System.Void Hast::InternalInvocationProxy().System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment) start
    -- Signal connections for Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0 (#0):
    \Unum::.ctor(UnumEnvironment).0._Started\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment)._Started.0\;
    \Unum::.ctor(UnumEnvironment).0.this.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment).this.parameter.Out.0\;
    \Unum::.ctor(UnumEnvironment).0.environment.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment).environment.parameter.Out.0\;
    \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment)._Finished.0\ <= \Unum::.ctor(UnumEnvironment).0._Finished\;
    \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment).this.parameter.In.0\ <= \Unum::.ctor(UnumEnvironment).0.this.parameter.Out\;
    \Unum::AddExactUnums(Unum,Unum).0.Unum::.ctor(UnumEnvironment).environment.parameter.In.0\ <= \Unum::.ctor(UnumEnvironment).0.environment.parameter.Out\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Lombiq.Unum.Unum::.ctor(Lombiq.Unum.UnumEnvironment) end


    -- System.Void Hast::InternalInvocationProxy().System.UInt16 Lombiq.Unum.Unum::get_FractionSizeMax() start
    -- Signal connections for Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0 (#0):
    \Unum::get_FractionSizeMax().0._Started\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Started.0\;
    \Unum::get_FractionSizeMax().0.this.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax().this.parameter.Out.0\;
    \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax()._Finished.0\ <= \Unum::get_FractionSizeMax().0._Finished\;
    \Unum::AddExactUnums(Unum,Unum).0.Unum::get_FractionSizeMax().return.0\ <= \Unum::get_FractionSizeMax().0.return\;
    -- System.Void Hast::InternalInvocationProxy().System.UInt16 Lombiq.Unum.Unum::get_FractionSizeMax() end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::AddAlignedFractions(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean) start
    -- Signal connections for Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0 (#0):
    \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._Started\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean)._Started.0\;
    \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.left.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean).left.parameter.Out.0\;
    \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.right.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean).right.parameter.Out.0\;
    \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.signBitsMatch.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean).signBitsMatch.parameter.Out.0\;
    \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean)._Finished.0\ <= \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0._Finished\;
    \Unum::AddExactUnums(Unum,Unum).0.Unum::AddAlignedFractions(BitMask,BitMask,Boolean).return.0\ <= \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.return\;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::AddAlignedFractions(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean) end


    -- System.Void Hast::InternalInvocationProxy().System.Boolean Lombiq.Unum.BitMask::op_GreaterThanOrEqual(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask) start
    -- Signal connections for Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0 (#0):
    \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._Started\ <= \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_GreaterThanOrEqual(BitMask,BitMask)._Started.0\;
    \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.left.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_GreaterThanOrEqual(BitMask,BitMask).left.parameter.Out.0\;
    \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.right.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_GreaterThanOrEqual(BitMask,BitMask).right.parameter.Out.0\;
    \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_GreaterThanOrEqual(BitMask,BitMask)._Finished.0\ <= \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0._Finished\;
    \Unum::AddExactUnums(Unum,Unum).0.BitMask::op_GreaterThanOrEqual(BitMask,BitMask).return.0\ <= \BitMask::op_GreaterThanOrEqual(BitMask,BitMask).0.return\;
    -- System.Void Hast::InternalInvocationProxy().System.Boolean Lombiq.Unum.BitMask::op_GreaterThanOrEqual(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask) end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentValueToExponentBits(System.Int32,System.Byte) start
    -- Signal connections for Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0 (#0):
    \Unum::ExponentValueToExponentBits(Int32,Byte).0._Started\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueToExponentBits(Int32,Byte)._Started.0\;
    \Unum::ExponentValueToExponentBits(Int32,Byte).0.value.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueToExponentBits(Int32,Byte).value.parameter.Out.0\;
    \Unum::ExponentValueToExponentBits(Int32,Byte).0.size.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueToExponentBits(Int32,Byte).size.parameter.Out.0\;
    \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueToExponentBits(Int32,Byte)._Finished.0\ <= \Unum::ExponentValueToExponentBits(Int32,Byte).0._Finished\;
    \Unum::AddExactUnums(Unum,Unum).0.Unum::ExponentValueToExponentBits(Int32,Byte).return.0\ <= \Unum::ExponentValueToExponentBits(Int32,Byte).0.return\;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.Unum::ExponentValueToExponentBits(System.Int32,System.Byte) end


    -- System.Void Hast::InternalInvocationProxy().System.Boolean Lombiq.Unum.Unum::IsExact() start
    -- Signal connections for Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0 (#0):
    \Unum::IsExact().0._Started\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::IsExact()._Started.0\;
    \Unum::IsExact().0.this.parameter.In\ <= \Unum::AddExactUnums(Unum,Unum).0.Unum::IsExact().this.parameter.Out.0\;
    \Unum::AddExactUnums(Unum,Unum).0.Unum::IsExact()._Finished.0\ <= \Unum::IsExact().0._Finished\;
    \Unum::AddExactUnums(Unum,Unum).0.Unum::IsExact().return.0\ <= \Unum::IsExact().0.return\;
    -- System.Void Hast::InternalInvocationProxy().System.Boolean Lombiq.Unum.Unum::IsExact() end


    -- System.Void Hast::InternalInvocationProxy().System.Boolean Lombiq.Unum.BitMask::op_GreaterThan(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask) start
    -- Signal connections for Lombiq.Unum.BitMask Lombiq.Unum.Unum::AddAlignedFractions(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask,System.Boolean).0 (#0):
    \BitMask::op_GreaterThan(BitMask,BitMask).0._Started\ <= \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_GreaterThan(BitMask,BitMask)._Started.0\;
    \BitMask::op_GreaterThan(BitMask,BitMask).0.left.parameter.In\ <= \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_GreaterThan(BitMask,BitMask).left.parameter.Out.0\;
    \BitMask::op_GreaterThan(BitMask,BitMask).0.right.parameter.In\ <= \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_GreaterThan(BitMask,BitMask).right.parameter.Out.0\;
    \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_GreaterThan(BitMask,BitMask)._Finished.0\ <= \BitMask::op_GreaterThan(BitMask,BitMask).0._Finished\;
    \Unum::AddAlignedFractions(BitMask,BitMask,Boolean).0.BitMask::op_GreaterThan(BitMask,BitMask).return.0\ <= \BitMask::op_GreaterThan(BitMask,BitMask).0.return\;
    -- System.Void Hast::InternalInvocationProxy().System.Boolean Lombiq.Unum.BitMask::op_GreaterThan(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask) end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum) start
    -- Signal connections for Lombiq.Unum.Unum Lombiq.Unum.Unum::op_Addition(Lombiq.Unum.Unum,Lombiq.Unum.Unum).0 (#0):
    \Unum::AddExactUnums(Unum,Unum).0._Started\ <= \Unum::op_Addition(Unum,Unum).0.Unum::AddExactUnums(Unum,Unum)._Started.0\;
    \Unum::AddExactUnums(Unum,Unum).0.left.parameter.In\ <= \Unum::op_Addition(Unum,Unum).0.Unum::AddExactUnums(Unum,Unum).left.parameter.Out.0\;
    \Unum::AddExactUnums(Unum,Unum).0.right.parameter.In\ <= \Unum::op_Addition(Unum,Unum).0.Unum::AddExactUnums(Unum,Unum).right.parameter.Out.0\;
    \Unum::op_Addition(Unum,Unum).0.Unum::AddExactUnums(Unum,Unum)._Finished.0\ <= \Unum::AddExactUnums(Unum,Unum).0._Finished\;
    \Unum::op_Addition(Unum,Unum).0.Unum::AddExactUnums(Unum,Unum).return.0\ <= \Unum::AddExactUnums(Unum,Unum).0.return\;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.Unum Lombiq.Unum.Unum::AddExactUnums(Lombiq.Unum.Unum,Lombiq.Unum.Unum) end


    -- System.Void Hast::InternalInvocationProxy().System.UInt16 Lombiq.Unum.UnumHelper::SegmentSizeSizeToSegmentSize(System.Byte) start
    -- Signal connections for System.Void Lombiq.Unum.UnumEnvironment::.ctor(System.Byte,System.Byte).0 (#0):
    \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._Started\ <= \UnumEnvironment::.ctor(Byte,Byte).0.UnumHelper::SegmentSizeSizeToSegmentSize(Byte)._Started.0\;
    \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0.segmentSizeSize.parameter.In\ <= \UnumEnvironment::.ctor(Byte,Byte).0.UnumHelper::SegmentSizeSizeToSegmentSize(Byte).segmentSizeSize.parameter.Out.0\;
    \UnumEnvironment::.ctor(Byte,Byte).0.UnumHelper::SegmentSizeSizeToSegmentSize(Byte)._Finished.0\ <= \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0._Finished\;
    \UnumEnvironment::.ctor(Byte,Byte).0.UnumHelper::SegmentSizeSizeToSegmentSize(Byte).return.0\ <= \UnumHelper::SegmentSizeSizeToSegmentSize(Byte).0.return\;
    -- System.Void Hast::InternalInvocationProxy().System.UInt16 Lombiq.Unum.UnumHelper::SegmentSizeSizeToSegmentSize(System.Byte) end


    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseOr(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask) start
    -- Signal connections for System.Void Lombiq.Unum.UnumEnvironment::.ctor(System.Byte,System.Byte).0 (#0):
    \BitMask::op_BitwiseOr(BitMask,BitMask).0._Started\ <= \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_BitwiseOr(BitMask,BitMask)._Started.0\;
    \BitMask::op_BitwiseOr(BitMask,BitMask).0.left.parameter.In\ <= \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_BitwiseOr(BitMask,BitMask).left.parameter.Out.0\;
    \BitMask::op_BitwiseOr(BitMask,BitMask).0.right.parameter.In\ <= \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_BitwiseOr(BitMask,BitMask).right.parameter.Out.0\;
    \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_BitwiseOr(BitMask,BitMask)._Finished.0\ <= \BitMask::op_BitwiseOr(BitMask,BitMask).0._Finished\;
    \UnumEnvironment::.ctor(Byte,Byte).0.BitMask::op_BitwiseOr(BitMask,BitMask).return.0\ <= \BitMask::op_BitwiseOr(BitMask,BitMask).0.return\;
    -- System.Void Hast::InternalInvocationProxy().Lombiq.Unum.BitMask Lombiq.Unum.BitMask::op_BitwiseOr(Lombiq.Unum.BitMask,Lombiq.Unum.BitMask) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.UnumCalculator::CalculateSumOfPowersofTwo(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._Started\ <= \Hast::ExternalInvocationProxy().UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory)._Started.0\;
    \Hast::ExternalInvocationProxy().UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory)._Finished.0\ <= \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.Samples.SampleAssembly.UnumCalculator::CalculateSumOfPowersofTwo(Hast.Transformer.Abstractions.SimpleMemory.SimpleMemory) end


    -- System.Void Hast::SimpleMemoryOperationProxy() start
    \CellIndex\ <= to_integer(\UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.SimpleMemory.CellIndex\) when \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.SimpleMemory.ReadEnable\ or \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.SimpleMemory.WriteEnable\ else 0;
    \DataOut\ <= \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.SimpleMemory.DataOut\ when \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.SimpleMemory.WriteEnable\ else "00000000000000000000000000000000";
    \ReadEnable\ <= \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.SimpleMemory.ReadEnable\;
    \WriteEnable\ <= \UnumCalculator::CalculateSumOfPowersofTwo(SimpleMemory).0.SimpleMemory.WriteEnable\;
    -- System.Void Hast::SimpleMemoryOperationProxy() end

end Imp;
