
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package TypeConversion is
	function Truncate(input: unsigned; size: natural) return unsigned;
	function Truncate(input: signed; size: natural) return signed;
end TypeConversion;
		
package body TypeConversion is

	function Truncate(input: unsigned; size: natural) return unsigned is
	begin
		return input(size - 1 downto 0);
	end Truncate;
	
	function Truncate(input: signed; size: natural) return signed is
	begin
		return input(size - 1 downto 0);
	end Truncate;

end TypeConversion;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.TypeConversion.all;

entity Hast_IP is 
    port(
        \MemberId\: In integer;
        \Reset\: In std_logic;
        \Started\: In boolean;
        \Finished\: Out boolean;
        \Clock\: In std_logic
    );
    -- (Hast_IP ID removed for approval testing.)
    -- (Date and time removed for approval testing.)
    -- Generated by Hastlayer - hastlayer.com
end Hast_IP;

architecture Imp of Hast_IP is 
    -- This IP was generated by Hastlayer from .NET code to mimic the original logic. Note the following:
    -- * For each member (methods, functions) in .NET a state machine was generated. Each state machine's name corresponds to 
    --   the original member's name.
    -- * Inputs and outputs are passed between state machines as shared objects.
    -- * There are operations that take multiple clock cycles like interacting with the memory and long-running arithmetic operations 
    --   (modulo, division, multiplication). These are awaited in subsequent states but be aware that some states can take more 
    --   than one clock cycle to produce their output.
    -- * The ExternalInvocationProxy process dispatches invocations that were started from the outside to the state machines.
    -- * The InternalInvocationProxy processes dispatch invocations between state machines.

    -- Custom inter-dependent type declarations start
    type \signed32_Array\ is array (integer range <>) of signed(31 downto 0);
    type \unsigned32_Array\ is array (integer range <>) of unsigned(31 downto 0);
    type \boolean_Array\ is array (integer range <>) of boolean;
    type \Hast.TestInputs.Various.ArrayUsingCases/ArrayHolder\ is record 
        \IsNull\: boolean;
        \Array\: \signed32_Array\(0 to 4);
    end record;
    type \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\ is record 
        \IsNull\: boolean;
        \ArrayLength\: unsigned(31 downto 0);
        \ArrayLengthCopy\: unsigned(31 downto 0);
        \NonSubstitutableArrayLengthCopy\: unsigned(31 downto 0);
        \Array\: \unsigned32_Array\(0 to 4);
    end record;
    type \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder2\ is record 
        \IsNull\: boolean;
        \ArrayLength\: unsigned(31 downto 0);
    end record;
    type \Hast.TestInputs.Various.ObjectUsingCases/MyClass\ is record 
        \IsNull\: boolean;
        \MyProperty\: signed(31 downto 0);
    end record;
    type \Hast.TestInputs.Various.ParallelCases/Calculator\ is record 
        \IsNull\: boolean;
        \Number\: unsigned(31 downto 0);
    end record;
    -- Custom inter-dependent type declarations end


    -- System.Void Hast.TestInputs.ClassStructure1.RootClass::VirtualMethod(System.Int32).0 declarations start
    -- State machine states:
    type \RootClass::VirtualMethod(Int32).0._States\ is (
        \RootClass::VirtualMethod(Int32).0._State_0\, 
        \RootClass::VirtualMethod(Int32).0._State_1\, 
        \RootClass::VirtualMethod(Int32).0._State_2\);
    -- Signals:
    Signal \RootClass::VirtualMethod(Int32).0._Finished\: boolean := false;
    Signal \RootClass::VirtualMethod(Int32).0._Started\: boolean := false;
    Signal \RootClass::VirtualMethod(Int32).0.input.parameter.In\: signed(31 downto 0) := to_signed(0, 32);
    -- System.Void Hast.TestInputs.ClassStructure1.RootClass::VirtualMethod(System.Int32).0 declarations end


    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0 declarations start
    -- State machine states:
    type \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._States\ is (
        \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._State_0\, 
        \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._State_1\, 
        \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._State_2\, 
        \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._State_3\);
    -- Signals:
    Signal \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._Finished\: boolean := false;
    Signal \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0.ComplexTypeHierarchy::PrivateMethod()._Started.0\: boolean := false;
    Signal \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._Started\: boolean := false;
    Signal \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0.ComplexTypeHierarchy::PrivateMethod()._Finished.0\: boolean := false;
    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0 declarations end


    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Interface1Method2().0 declarations start
    -- State machine states:
    type \ComplexTypeHierarchy::Interface1Method2().0._States\ is (
        \ComplexTypeHierarchy::Interface1Method2().0._State_0\, 
        \ComplexTypeHierarchy::Interface1Method2().0._State_1\, 
        \ComplexTypeHierarchy::Interface1Method2().0._State_2\, 
        \ComplexTypeHierarchy::Interface1Method2().0._State_3\, 
        \ComplexTypeHierarchy::Interface1Method2().0._State_4\);
    -- Signals:
    Signal \ComplexTypeHierarchy::Interface1Method2().0._Finished\: boolean := false;
    Signal \ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::PrivateMethod()._Started.0\: boolean := false;
    Signal \ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::StaticMethod()._Started.0\: boolean := false;
    Signal \ComplexTypeHierarchy::Interface1Method2().0._Started\: boolean := false;
    Signal \ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::PrivateMethod()._Finished.0\: boolean := false;
    Signal \ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::StaticMethod()._Finished.0\: boolean := false;
    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Interface1Method2().0 declarations end


    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Interface2Method1().0 declarations start
    -- State machine states:
    type \ComplexTypeHierarchy::Interface2Method1().0._States\ is (
        \ComplexTypeHierarchy::Interface2Method1().0._State_0\, 
        \ComplexTypeHierarchy::Interface2Method1().0._State_1\, 
        \ComplexTypeHierarchy::Interface2Method1().0._State_2\, 
        \ComplexTypeHierarchy::Interface2Method1().0._State_3\);
    -- Signals:
    Signal \ComplexTypeHierarchy::Interface2Method1().0._Finished\: boolean := false;
    Signal \ComplexTypeHierarchy::Interface2Method1().0.ComplexTypeHierarchy::BaseInterfaceMethod2()._Started.0\: boolean := false;
    Signal \ComplexTypeHierarchy::Interface2Method1().0._Started\: boolean := false;
    Signal \ComplexTypeHierarchy::Interface2Method1().0.ComplexTypeHierarchy::BaseInterfaceMethod2()._Finished.0\: boolean := false;
    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Interface2Method1().0 declarations end


    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0 declarations start
    -- State machine states:
    type \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._States\ is (
        \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._State_0\, 
        \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._State_1\, 
        \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._State_2\);
    -- Signals:
    Signal \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._Finished\: boolean := false;
    Signal \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._Started\: boolean := false;
    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0 declarations end


    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::BaseInterfaceMethod2().0 declarations start
    -- State machine states:
    type \ComplexTypeHierarchy::BaseInterfaceMethod2().0._States\ is (
        \ComplexTypeHierarchy::BaseInterfaceMethod2().0._State_0\, 
        \ComplexTypeHierarchy::BaseInterfaceMethod2().0._State_1\, 
        \ComplexTypeHierarchy::BaseInterfaceMethod2().0._State_2\, 
        \ComplexTypeHierarchy::BaseInterfaceMethod2().0._State_3\);
    -- Signals:
    Signal \ComplexTypeHierarchy::BaseInterfaceMethod2().0._Finished\: boolean := false;
    Signal \ComplexTypeHierarchy::BaseInterfaceMethod2().0.ComplexTypeHierarchy::StaticMethod()._Started.0\: boolean := false;
    Signal \ComplexTypeHierarchy::BaseInterfaceMethod2().0._Started\: boolean := false;
    Signal \ComplexTypeHierarchy::BaseInterfaceMethod2().0.ComplexTypeHierarchy::StaticMethod()._Finished.0\: boolean := false;
    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::BaseInterfaceMethod2().0 declarations end


    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0 declarations start
    -- State machine states:
    type \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._States\ is (
        \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._State_0\, 
        \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._State_1\, 
        \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._State_2\, 
        \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._State_3\);
    -- Signals:
    Signal \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._Finished\: boolean := false;
    Signal \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0.ComplexTypeHierarchy::PrivateMethod()._Started.0\: boolean := false;
    Signal \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._Started\: boolean := false;
    Signal \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0.ComplexTypeHierarchy::PrivateMethod()._Finished.0\: boolean := false;
    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0 declarations end


    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::PrivateMethod().0 declarations start
    -- State machine states:
    type \ComplexTypeHierarchy::PrivateMethod().0._States\ is (
        \ComplexTypeHierarchy::PrivateMethod().0._State_0\, 
        \ComplexTypeHierarchy::PrivateMethod().0._State_1\, 
        \ComplexTypeHierarchy::PrivateMethod().0._State_2\, 
        \ComplexTypeHierarchy::PrivateMethod().0._State_3\);
    -- Signals:
    Signal \ComplexTypeHierarchy::PrivateMethod().0._Finished\: boolean := false;
    Signal \ComplexTypeHierarchy::PrivateMethod().0.ComplexTypeHierarchy::StaticMethod()._Started.0\: boolean := false;
    Signal \ComplexTypeHierarchy::PrivateMethod().0._Started\: boolean := false;
    Signal \ComplexTypeHierarchy::PrivateMethod().0.ComplexTypeHierarchy::StaticMethod()._Finished.0\: boolean := false;
    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::PrivateMethod().0 declarations end


    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::StaticMethod().0 declarations start
    -- State machine states:
    type \ComplexTypeHierarchy::StaticMethod().0._States\ is (
        \ComplexTypeHierarchy::StaticMethod().0._State_0\, 
        \ComplexTypeHierarchy::StaticMethod().0._State_1\, 
        \ComplexTypeHierarchy::StaticMethod().0._State_2\);
    -- Signals:
    Signal \ComplexTypeHierarchy::StaticMethod().0._Finished\: boolean := false;
    Signal \ComplexTypeHierarchy::StaticMethod().0._Started\: boolean := false;
    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::StaticMethod().0 declarations end


    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.StaticClass::StaticMethod().0 declarations start
    -- State machine states:
    type \StaticClass::StaticMethod().0._States\ is (
        \StaticClass::StaticMethod().0._State_0\, 
        \StaticClass::StaticMethod().0._State_1\, 
        \StaticClass::StaticMethod().0._State_2\);
    -- Signals:
    Signal \StaticClass::StaticMethod().0._Finished\: boolean := false;
    Signal \StaticClass::StaticMethod().0._Started\: boolean := false;
    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.StaticClass::StaticMethod().0 declarations end


    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.UnusedDeclarations::UnusedMethod().0 declarations start
    -- State machine states:
    type \UnusedDeclarations::UnusedMethod().0._States\ is (
        \UnusedDeclarations::UnusedMethod().0._State_0\, 
        \UnusedDeclarations::UnusedMethod().0._State_1\, 
        \UnusedDeclarations::UnusedMethod().0._State_2\);
    -- Signals:
    Signal \UnusedDeclarations::UnusedMethod().0._Finished\: boolean := false;
    Signal \UnusedDeclarations::UnusedMethod().0._Started\: boolean := false;
    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.UnusedDeclarations::UnusedMethod().0 declarations end


    -- System.Void Hast.TestInputs.ClassStructure2.StaticReference::StaticClassUsingMethod().0 declarations start
    -- State machine states:
    type \StaticReference::StaticClassUsingMethod().0._States\ is (
        \StaticReference::StaticClassUsingMethod().0._State_0\, 
        \StaticReference::StaticClassUsingMethod().0._State_1\, 
        \StaticReference::StaticClassUsingMethod().0._State_2\, 
        \StaticReference::StaticClassUsingMethod().0._State_3\);
    -- Signals:
    Signal \StaticReference::StaticClassUsingMethod().0._Finished\: boolean := false;
    Signal \StaticReference::StaticClassUsingMethod().0.StaticClass::StaticMethod()._Started.0\: boolean := false;
    Signal \StaticReference::StaticClassUsingMethod().0._Started\: boolean := false;
    Signal \StaticReference::StaticClassUsingMethod().0.StaticClass::StaticMethod()._Finished.0\: boolean := false;
    -- System.Void Hast.TestInputs.ClassStructure2.StaticReference::StaticClassUsingMethod().0 declarations end


    -- System.Void Hast.TestInputs.Various.ArrayUsingCases/ArrayHolder::.ctor(System.Int32[]).0 declarations start
    -- State machine states:
    type \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._States\ is (
        \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._State_0\, 
        \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._State_1\, 
        \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._State_2\);
    -- Signals:
    Signal \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._Finished\: boolean := false;
    Signal \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0.this.parameter.Out\: \Hast.TestInputs.Various.ArrayUsingCases/ArrayHolder\;
    Signal \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0.array.parameter.Out\: \signed32_Array\(0 to 4) := (others => to_signed(0, 32));
    Signal \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._Started\: boolean := false;
    Signal \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0.this.parameter.In\: \Hast.TestInputs.Various.ArrayUsingCases/ArrayHolder\;
    Signal \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0.array.parameter.In\: \signed32_Array\(0 to 4) := (others => to_signed(0, 32));
    -- System.Void Hast.TestInputs.Various.ArrayUsingCases/ArrayHolder::.ctor(System.Int32[]).0 declarations end


    -- System.Void Hast.TestInputs.Various.ArrayUsingCases::PassArrayToConstructor().0 declarations start
    -- State machine states:
    type \ArrayUsingCases::PassArrayToConstructor().0._States\ is (
        \ArrayUsingCases::PassArrayToConstructor().0._State_0\, 
        \ArrayUsingCases::PassArrayToConstructor().0._State_1\, 
        \ArrayUsingCases::PassArrayToConstructor().0._State_2\, 
        \ArrayUsingCases::PassArrayToConstructor().0._State_3\);
    -- Signals:
    Signal \ArrayUsingCases::PassArrayToConstructor().0._Finished\: boolean := false;
    Signal \ArrayUsingCases::PassArrayToConstructor().0.ArrayUsingCases/ArrayHolder::.ctor(Int32[]).this.parameter.Out.0\: \Hast.TestInputs.Various.ArrayUsingCases/ArrayHolder\;
    Signal \ArrayUsingCases::PassArrayToConstructor().0.ArrayUsingCases/ArrayHolder::.ctor(Int32[]).array.parameter.Out.0\: \signed32_Array\(0 to 4) := (others => to_signed(0, 32));
    Signal \ArrayUsingCases::PassArrayToConstructor().0.ArrayUsingCases/ArrayHolder::.ctor(Int32[])._Started.0\: boolean := false;
    Signal \ArrayUsingCases::PassArrayToConstructor().0._Started\: boolean := false;
    Signal \ArrayUsingCases::PassArrayToConstructor().0.ArrayUsingCases/ArrayHolder::.ctor(Int32[]).this.parameter.In.0\: \Hast.TestInputs.Various.ArrayUsingCases/ArrayHolder\;
    Signal \ArrayUsingCases::PassArrayToConstructor().0.ArrayUsingCases/ArrayHolder::.ctor(Int32[]).array.parameter.In.0\: \signed32_Array\(0 to 4) := (others => to_signed(0, 32));
    Signal \ArrayUsingCases::PassArrayToConstructor().0.ArrayUsingCases/ArrayHolder::.ctor(Int32[])._Finished.0\: boolean := false;
    -- System.Void Hast.TestInputs.Various.ArrayUsingCases::PassArrayToConstructor().0 declarations end


    -- System.Void Hast.TestInputs.Various.ArrayUsingCases::PassArrayFromMethod().0 declarations start
    -- State machine states:
    type \ArrayUsingCases::PassArrayFromMethod().0._States\ is (
        \ArrayUsingCases::PassArrayFromMethod().0._State_0\, 
        \ArrayUsingCases::PassArrayFromMethod().0._State_1\, 
        \ArrayUsingCases::PassArrayFromMethod().0._State_2\, 
        \ArrayUsingCases::PassArrayFromMethod().0._State_3\);
    -- Signals:
    Signal \ArrayUsingCases::PassArrayFromMethod().0._Finished\: boolean := false;
    Signal \ArrayUsingCases::PassArrayFromMethod().0.ArrayUsingCases::ArrayProducingMethod(Int32).arrayLength.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \ArrayUsingCases::PassArrayFromMethod().0.ArrayUsingCases::ArrayProducingMethod(Int32)._Started.0\: boolean := false;
    Signal \ArrayUsingCases::PassArrayFromMethod().0._Started\: boolean := false;
    Signal \ArrayUsingCases::PassArrayFromMethod().0.ArrayUsingCases::ArrayProducingMethod(Int32)._Finished.0\: boolean := false;
    Signal \ArrayUsingCases::PassArrayFromMethod().0.ArrayUsingCases::ArrayProducingMethod(Int32).return.0\: \signed32_Array\(0 to 4) := (others => to_signed(0, 32));
    -- System.Void Hast.TestInputs.Various.ArrayUsingCases::PassArrayFromMethod().0 declarations end


    -- System.Int32[] Hast.TestInputs.Various.ArrayUsingCases::ArrayProducingMethod(System.Int32).0 declarations start
    -- State machine states:
    type \ArrayUsingCases::ArrayProducingMethod(Int32).0._States\ is (
        \ArrayUsingCases::ArrayProducingMethod(Int32).0._State_0\, 
        \ArrayUsingCases::ArrayProducingMethod(Int32).0._State_1\, 
        \ArrayUsingCases::ArrayProducingMethod(Int32).0._State_2\);
    -- Signals:
    Signal \ArrayUsingCases::ArrayProducingMethod(Int32).0._Finished\: boolean := false;
    Signal \ArrayUsingCases::ArrayProducingMethod(Int32).0.return\: \signed32_Array\(0 to 4) := (others => to_signed(0, 32));
    Signal \ArrayUsingCases::ArrayProducingMethod(Int32).0._Started\: boolean := false;
    Signal \ArrayUsingCases::ArrayProducingMethod(Int32).0.arrayLength.parameter.In\: signed(31 downto 0) := to_signed(0, 32);
    -- System.Int32[] Hast.TestInputs.Various.ArrayUsingCases::ArrayProducingMethod(System.Int32).0 declarations end


    -- System.Void Hast.TestInputs.Various.CastingCases::NumberCasting(System.Int16,System.Int16).0 declarations start
    -- State machine states:
    type \CastingCases::NumberCasting(Int16,Int16).0._States\ is (
        \CastingCases::NumberCasting(Int16,Int16).0._State_0\, 
        \CastingCases::NumberCasting(Int16,Int16).0._State_1\, 
        \CastingCases::NumberCasting(Int16,Int16).0._State_2\);
    -- Signals:
    Signal \CastingCases::NumberCasting(Int16,Int16).0._Finished\: boolean := false;
    Signal \CastingCases::NumberCasting(Int16,Int16).0._Started\: boolean := false;
    Signal \CastingCases::NumberCasting(Int16,Int16).0.a.parameter.In\: signed(15 downto 0) := to_signed(0, 16);
    Signal \CastingCases::NumberCasting(Int16,Int16).0.b.parameter.In\: signed(15 downto 0) := to_signed(0, 16);
    -- System.Void Hast.TestInputs.Various.CastingCases::NumberCasting(System.Int16,System.Int16).0 declarations end


    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32[]).0 declarations start
    -- State machine states:
    type \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._States\ is (
        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._State_0\, 
        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._State_1\, 
        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._State_2\);
    -- Signals:
    Signal \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._Finished\: boolean := false;
    Signal \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.this.parameter.Out\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
    Signal \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.array.parameter.Out\: \unsigned32_Array\(0 to 4) := (others => to_unsigned(0, 32));
    Signal \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._Started\: boolean := false;
    Signal \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.this.parameter.In\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
    Signal \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.array.parameter.In\: \unsigned32_Array\(0 to 4) := (others => to_unsigned(0, 32));
    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32[]).0 declarations end


    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32).0 declarations start
    -- State machine states:
    type \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._States\ is (
        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._State_0\, 
        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._State_1\, 
        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._State_2\);
    -- Signals:
    Signal \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._Finished\: boolean := false;
    Signal \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0.this.parameter.Out\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
    Signal \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._Started\: boolean := false;
    Signal \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0.this.parameter.In\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
    Signal \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0.size.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32).0 declarations end


    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1).0 declarations start
    -- State machine states:
    type \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._States\ is (
        \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._State_0\, 
        \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._State_1\, 
        \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._State_2\, 
        \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._State_3\);
    -- Signals:
    Signal \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._Finished\: boolean := false;
    Signal \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.this.parameter.Out\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
    Signal \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.previous.parameter.Out\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
    Signal \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).this.parameter.Out.0\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
    Signal \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).array.parameter.Out.0\: \unsigned32_Array\(0 to 4) := (others => to_unsigned(0, 32));
    Signal \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Started.0\: boolean := false;
    Signal \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._Started\: boolean := false;
    Signal \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.this.parameter.In\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
    Signal \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.previous.parameter.In\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
    Signal \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).this.parameter.In.0\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
    Signal \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).array.parameter.In.0\: \unsigned32_Array\(0 to 4) := (others => to_unsigned(0, 32));
    Signal \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Finished.0\: boolean := false;
    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1).0 declarations end


    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder2::.ctor(System.UInt32).0 declarations start
    -- State machine states:
    type \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._States\ is (
        \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_0\, 
        \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_1\, 
        \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_2\, 
        \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_3\, 
        \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_4\, 
        \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_5\, 
        \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_6\, 
        \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_7\);
    -- Signals:
    Signal \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._Finished\: boolean := false;
    Signal \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.this.parameter.Out\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder2\;
    Signal \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._Started\: boolean := false;
    Signal \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.this.parameter.In\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder2\;
    Signal \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.size.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder2::.ctor(System.UInt32).0 declarations end


    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases::ConstantValuedVariables(System.Int32).0 declarations start
    -- State machine states:
    type \ConstantsUsingCases::ConstantValuedVariables(Int32).0._States\ is (
        \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_0\, 
        \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_1\, 
        \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_2\, 
        \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_3\, 
        \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_4\);
    -- Signals:
    Signal \ConstantsUsingCases::ConstantValuedVariables(Int32).0._Finished\: boolean := false;
    Signal \ConstantsUsingCases::ConstantValuedVariables(Int32).0._Started\: boolean := false;
    Signal \ConstantsUsingCases::ConstantValuedVariables(Int32).0.input.parameter.In\: signed(31 downto 0) := to_signed(0, 32);
    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases::ConstantValuedVariables(System.Int32).0 declarations end


    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases::ConstantPassingToMethod(System.Int32).0 declarations start
    -- State machine states:
    type \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._States\ is (
        \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._State_0\, 
        \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._State_1\, 
        \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._State_2\, 
        \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._State_3\);
    -- Signals:
    Signal \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._Finished\: boolean := false;
    Signal \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).input1.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).input2.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.ConstantsUsingCases::ConstantUsingMethod(Int32,Int32)._Started.0\: boolean := false;
    Signal \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._Started\: boolean := false;
    Signal \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.input.parameter.In\: signed(31 downto 0) := to_signed(0, 32);
    Signal \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.ConstantsUsingCases::ConstantUsingMethod(Int32,Int32)._Finished.0\: boolean := false;
    Signal \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).return.0\: signed(31 downto 0) := to_signed(0, 32);
    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases::ConstantPassingToMethod(System.Int32).0 declarations end


    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases::ConstantPassingToObject().0 declarations start
    -- State machine states:
    type \ConstantsUsingCases::ConstantPassingToObject().0._States\ is (
        \ConstantsUsingCases::ConstantPassingToObject().0._State_0\, 
        \ConstantsUsingCases::ConstantPassingToObject().0._State_1\, 
        \ConstantsUsingCases::ConstantPassingToObject().0._State_2\, 
        \ConstantsUsingCases::ConstantPassingToObject().0._State_3\, 
        \ConstantsUsingCases::ConstantPassingToObject().0._State_4\, 
        \ConstantsUsingCases::ConstantPassingToObject().0._State_5\, 
        \ConstantsUsingCases::ConstantPassingToObject().0._State_6\, 
        \ConstantsUsingCases::ConstantPassingToObject().0._State_7\, 
        \ConstantsUsingCases::ConstantPassingToObject().0._State_8\, 
        \ConstantsUsingCases::ConstantPassingToObject().0._State_9\, 
        \ConstantsUsingCases::ConstantPassingToObject().0._State_10\);
    -- Signals:
    Signal \ConstantsUsingCases::ConstantPassingToObject().0._Finished\: boolean := false;
    Signal \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).this.parameter.Out.0\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
    Signal \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).array.parameter.Out.0\: \unsigned32_Array\(0 to 4) := (others => to_unsigned(0, 32));
    Signal \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Started.0\: boolean := false;
    Signal \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).this.parameter.Out.0\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
    Signal \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).size.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32)._Started.0\: boolean := false;
    Signal \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).this.parameter.Out.0\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
    Signal \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).previous.parameter.Out.0\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
    Signal \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1)._Started.0\: boolean := false;
    Signal \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).this.parameter.Out.0\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder2\;
    Signal \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).size.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32)._Started.0\: boolean := false;
    Signal \ConstantsUsingCases::ConstantPassingToObject().0._Started\: boolean := false;
    Signal \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).this.parameter.In.0\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
    Signal \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).array.parameter.In.0\: \unsigned32_Array\(0 to 4) := (others => to_unsigned(0, 32));
    Signal \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Finished.0\: boolean := false;
    Signal \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).this.parameter.In.0\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
    Signal \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32)._Finished.0\: boolean := false;
    Signal \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).this.parameter.In.0\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
    Signal \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).previous.parameter.In.0\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
    Signal \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1)._Finished.0\: boolean := false;
    Signal \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).this.parameter.In.0\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder2\;
    Signal \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32)._Finished.0\: boolean := false;
    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases::ConstantPassingToObject().0 declarations end


    -- System.Int32 Hast.TestInputs.Various.ConstantsUsingCases::ConstantUsingMethod(System.Int32,System.Int32).0 declarations start
    -- State machine states:
    type \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._States\ is (
        \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._State_0\, 
        \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._State_1\, 
        \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._State_2\);
    -- Signals:
    Signal \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._Finished\: boolean := false;
    Signal \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0.return\: signed(31 downto 0) := to_signed(0, 32);
    Signal \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._Started\: boolean := false;
    Signal \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0.input1.parameter.In\: signed(31 downto 0) := to_signed(0, 32);
    Signal \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0.input2.parameter.In\: signed(31 downto 0) := to_signed(0, 32);
    -- System.Int32 Hast.TestInputs.Various.ConstantsUsingCases::ConstantUsingMethod(System.Int32,System.Int32).0 declarations end


    -- System.Void Hast.TestInputs.Various.LoopCases::BreakInLoop(System.Int32).0 declarations start
    -- State machine states:
    type \LoopCases::BreakInLoop(Int32).0._States\ is (
        \LoopCases::BreakInLoop(Int32).0._State_0\, 
        \LoopCases::BreakInLoop(Int32).0._State_1\, 
        \LoopCases::BreakInLoop(Int32).0._State_2\, 
        \LoopCases::BreakInLoop(Int32).0._State_3\, 
        \LoopCases::BreakInLoop(Int32).0._State_4\, 
        \LoopCases::BreakInLoop(Int32).0._State_5\, 
        \LoopCases::BreakInLoop(Int32).0._State_6\);
    -- Signals:
    Signal \LoopCases::BreakInLoop(Int32).0._Finished\: boolean := false;
    Signal \LoopCases::BreakInLoop(Int32).0._Started\: boolean := false;
    Signal \LoopCases::BreakInLoop(Int32).0.input.parameter.In\: signed(31 downto 0) := to_signed(0, 32);
    -- System.Void Hast.TestInputs.Various.LoopCases::BreakInLoop(System.Int32).0 declarations end


    -- System.Void Hast.TestInputs.Various.LoopCases::BreakInLoopInLoop(System.Int32).0 declarations start
    -- State machine states:
    type \LoopCases::BreakInLoopInLoop(Int32).0._States\ is (
        \LoopCases::BreakInLoopInLoop(Int32).0._State_0\, 
        \LoopCases::BreakInLoopInLoop(Int32).0._State_1\, 
        \LoopCases::BreakInLoopInLoop(Int32).0._State_2\, 
        \LoopCases::BreakInLoopInLoop(Int32).0._State_3\, 
        \LoopCases::BreakInLoopInLoop(Int32).0._State_4\, 
        \LoopCases::BreakInLoopInLoop(Int32).0._State_5\, 
        \LoopCases::BreakInLoopInLoop(Int32).0._State_6\, 
        \LoopCases::BreakInLoopInLoop(Int32).0._State_7\, 
        \LoopCases::BreakInLoopInLoop(Int32).0._State_8\);
    -- Signals:
    Signal \LoopCases::BreakInLoopInLoop(Int32).0._Finished\: boolean := false;
    Signal \LoopCases::BreakInLoopInLoop(Int32).0._Started\: boolean := false;
    Signal \LoopCases::BreakInLoopInLoop(Int32).0.input.parameter.In\: signed(31 downto 0) := to_signed(0, 32);
    -- System.Void Hast.TestInputs.Various.LoopCases::BreakInLoopInLoop(System.Int32).0 declarations end


    -- System.Void Hast.TestInputs.Various.ObjectUsingCases::NullUsage().0 declarations start
    -- State machine states:
    type \ObjectUsingCases::NullUsage().0._States\ is (
        \ObjectUsingCases::NullUsage().0._State_0\, 
        \ObjectUsingCases::NullUsage().0._State_1\, 
        \ObjectUsingCases::NullUsage().0._State_2\, 
        \ObjectUsingCases::NullUsage().0._State_3\, 
        \ObjectUsingCases::NullUsage().0._State_4\, 
        \ObjectUsingCases::NullUsage().0._State_5\, 
        \ObjectUsingCases::NullUsage().0._State_6\);
    -- Signals:
    Signal \ObjectUsingCases::NullUsage().0._Finished\: boolean := false;
    Signal \ObjectUsingCases::NullUsage().0._Started\: boolean := false;
    -- System.Void Hast.TestInputs.Various.ObjectUsingCases::NullUsage().0 declarations end


    -- System.Void Hast.TestInputs.Various.ObjectUsingCases::VoidReturn(System.Int32).0 declarations start
    -- State machine states:
    type \ObjectUsingCases::VoidReturn(Int32).0._States\ is (
        \ObjectUsingCases::VoidReturn(Int32).0._State_0\, 
        \ObjectUsingCases::VoidReturn(Int32).0._State_1\, 
        \ObjectUsingCases::VoidReturn(Int32).0._State_2\, 
        \ObjectUsingCases::VoidReturn(Int32).0._State_3\);
    -- Signals:
    Signal \ObjectUsingCases::VoidReturn(Int32).0._Finished\: boolean := false;
    Signal \ObjectUsingCases::VoidReturn(Int32).0.ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).myClass.parameter.Out.0\: \Hast.TestInputs.Various.ObjectUsingCases/MyClass\;
    Signal \ObjectUsingCases::VoidReturn(Int32).0.ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass)._Started.0\: boolean := false;
    Signal \ObjectUsingCases::VoidReturn(Int32).0._Started\: boolean := false;
    Signal \ObjectUsingCases::VoidReturn(Int32).0.input.parameter.In\: signed(31 downto 0) := to_signed(0, 32);
    Signal \ObjectUsingCases::VoidReturn(Int32).0.ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).myClass.parameter.In.0\: \Hast.TestInputs.Various.ObjectUsingCases/MyClass\;
    Signal \ObjectUsingCases::VoidReturn(Int32).0.ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass)._Finished.0\: boolean := false;
    -- System.Void Hast.TestInputs.Various.ObjectUsingCases::VoidReturn(System.Int32).0 declarations end


    -- System.Void Hast.TestInputs.Various.ObjectUsingCases::VoidMethod(Hast.TestInputs.Various.ObjectUsingCases/MyClass).0 declarations start
    -- State machine states:
    type \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._States\ is (
        \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_0\, 
        \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_1\, 
        \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_2\, 
        \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_3\, 
        \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_4\, 
        \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_5\, 
        \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_6\);
    -- Signals:
    Signal \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._Finished\: boolean := false;
    Signal \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.myClass.parameter.Out\: \Hast.TestInputs.Various.ObjectUsingCases/MyClass\;
    Signal \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._Started\: boolean := false;
    Signal \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.myClass.parameter.In\: \Hast.TestInputs.Various.ObjectUsingCases/MyClass\;
    -- System.Void Hast.TestInputs.Various.ObjectUsingCases::VoidMethod(Hast.TestInputs.Various.ObjectUsingCases/MyClass).0 declarations end


    -- System.Boolean Hast.TestInputs.Various.ParallelCases/Calculator::IsEven().0 declarations start
    -- State machine states:
    type \ParallelCases/Calculator::IsEven().0._States\ is (
        \ParallelCases/Calculator::IsEven().0._State_0\, 
        \ParallelCases/Calculator::IsEven().0._State_1\, 
        \ParallelCases/Calculator::IsEven().0._State_2\, 
        \ParallelCases/Calculator::IsEven().0._State_3\, 
        \ParallelCases/Calculator::IsEven().0._State_4\);
    -- Signals:
    Signal \ParallelCases/Calculator::IsEven().0._Finished\: boolean := false;
    Signal \ParallelCases/Calculator::IsEven().0.return\: boolean := false;
    Signal \ParallelCases/Calculator::IsEven().0.this.parameter.Out\: \Hast.TestInputs.Various.ParallelCases/Calculator\;
    Signal \ParallelCases/Calculator::IsEven().0._Started\: boolean := false;
    Signal \ParallelCases/Calculator::IsEven().0.this.parameter.In\: \Hast.TestInputs.Various.ParallelCases/Calculator\;
    -- System.Boolean Hast.TestInputs.Various.ParallelCases/Calculator::IsEven().0 declarations end


    -- System.Boolean Hast.TestInputs.Various.ParallelCases/Calculator::IsEven().1 declarations start
    -- State machine states:
    type \ParallelCases/Calculator::IsEven().1._States\ is (
        \ParallelCases/Calculator::IsEven().1._State_0\, 
        \ParallelCases/Calculator::IsEven().1._State_1\, 
        \ParallelCases/Calculator::IsEven().1._State_2\, 
        \ParallelCases/Calculator::IsEven().1._State_3\, 
        \ParallelCases/Calculator::IsEven().1._State_4\);
    -- Signals:
    Signal \ParallelCases/Calculator::IsEven().1._Finished\: boolean := false;
    Signal \ParallelCases/Calculator::IsEven().1.return\: boolean := false;
    Signal \ParallelCases/Calculator::IsEven().1.this.parameter.Out\: \Hast.TestInputs.Various.ParallelCases/Calculator\;
    Signal \ParallelCases/Calculator::IsEven().1._Started\: boolean := false;
    Signal \ParallelCases/Calculator::IsEven().1.this.parameter.In\: \Hast.TestInputs.Various.ParallelCases/Calculator\;
    -- System.Boolean Hast.TestInputs.Various.ParallelCases/Calculator::IsEven().1 declarations end


    -- System.Boolean Hast.TestInputs.Various.ParallelCases/Calculator::IsEven().2 declarations start
    -- State machine states:
    type \ParallelCases/Calculator::IsEven().2._States\ is (
        \ParallelCases/Calculator::IsEven().2._State_0\, 
        \ParallelCases/Calculator::IsEven().2._State_1\, 
        \ParallelCases/Calculator::IsEven().2._State_2\, 
        \ParallelCases/Calculator::IsEven().2._State_3\, 
        \ParallelCases/Calculator::IsEven().2._State_4\);
    -- Signals:
    Signal \ParallelCases/Calculator::IsEven().2._Finished\: boolean := false;
    Signal \ParallelCases/Calculator::IsEven().2.return\: boolean := false;
    Signal \ParallelCases/Calculator::IsEven().2.this.parameter.Out\: \Hast.TestInputs.Various.ParallelCases/Calculator\;
    Signal \ParallelCases/Calculator::IsEven().2._Started\: boolean := false;
    Signal \ParallelCases/Calculator::IsEven().2.this.parameter.In\: \Hast.TestInputs.Various.ParallelCases/Calculator\;
    -- System.Boolean Hast.TestInputs.Various.ParallelCases/Calculator::IsEven().2 declarations end


    -- System.UInt32 Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::input declarations start
    -- Shared (global) variables:
    shared Variable \System.UInt32 Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::input\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.UInt32 Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::input declarations end


    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(System.UInt32).0 declarations start
    -- State machine states:
    type \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._States\ is (
        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State_0\, 
        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State_1\, 
        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State_2\, 
        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State_3\, 
        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State_4\);
    -- Signals:
    Signal \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._Finished\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.return\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._Started\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.indexObject.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(System.UInt32).0 declarations end


    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(System.UInt32).1 declarations start
    -- State machine states:
    type \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._States\ is (
        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State_0\, 
        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State_1\, 
        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State_2\, 
        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State_3\, 
        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State_4\);
    -- Signals:
    Signal \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._Finished\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.return\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._Started\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.indexObject.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(System.UInt32).1 declarations end


    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(System.UInt32).2 declarations start
    -- State machine states:
    type \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._States\ is (
        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State_0\, 
        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State_1\, 
        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State_2\, 
        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State_3\, 
        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State_4\);
    -- Signals:
    Signal \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._Finished\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.return\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._Started\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.indexObject.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(System.UInt32).2 declarations end


    -- System.UInt32 Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::input declarations start
    -- Shared (global) variables:
    shared Variable \System.UInt32 Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::input\: unsigned(31 downto 0) := to_unsigned(0, 32);
    -- System.UInt32 Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::input declarations end


    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(System.UInt32).0 declarations start
    -- State machine states:
    type \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._States\ is (
        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._State_0\, 
        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._State_1\, 
        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._State_2\, 
        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._State_3\);
    -- Signals:
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._Finished\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.return\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.ParallelCases/Calculator::IsEven().this.parameter.Out.0\: \Hast.TestInputs.Various.ParallelCases/Calculator\;
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.ParallelCases/Calculator::IsEven()._Started.0\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._Started\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.indexObject.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.ParallelCases/Calculator::IsEven().this.parameter.In.0\: \Hast.TestInputs.Various.ParallelCases/Calculator\;
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.ParallelCases/Calculator::IsEven()._Finished.0\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.ParallelCases/Calculator::IsEven().return.0\: boolean := false;
    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(System.UInt32).0 declarations end


    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(System.UInt32).1 declarations start
    -- State machine states:
    type \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._States\ is (
        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._State_0\, 
        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._State_1\, 
        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._State_2\, 
        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._State_3\);
    -- Signals:
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._Finished\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.return\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.ParallelCases/Calculator::IsEven().this.parameter.Out.0\: \Hast.TestInputs.Various.ParallelCases/Calculator\;
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.ParallelCases/Calculator::IsEven()._Started.0\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._Started\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.indexObject.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.ParallelCases/Calculator::IsEven().this.parameter.In.0\: \Hast.TestInputs.Various.ParallelCases/Calculator\;
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.ParallelCases/Calculator::IsEven()._Finished.0\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.ParallelCases/Calculator::IsEven().return.0\: boolean := false;
    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(System.UInt32).1 declarations end


    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(System.UInt32).2 declarations start
    -- State machine states:
    type \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._States\ is (
        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._State_0\, 
        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._State_1\, 
        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._State_2\, 
        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._State_3\);
    -- Signals:
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._Finished\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.return\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.ParallelCases/Calculator::IsEven().this.parameter.Out.0\: \Hast.TestInputs.Various.ParallelCases/Calculator\;
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.ParallelCases/Calculator::IsEven()._Started.0\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._Started\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.indexObject.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.ParallelCases/Calculator::IsEven().this.parameter.In.0\: \Hast.TestInputs.Various.ParallelCases/Calculator\;
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.ParallelCases/Calculator::IsEven()._Finished.0\: boolean := false;
    Signal \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.ParallelCases/Calculator::IsEven().return.0\: boolean := false;
    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(System.UInt32).2 declarations end


    -- System.Void Hast.TestInputs.Various.ParallelCases::WhenAllWhenAnyAwaitedTasks(System.UInt32).0 declarations start
    -- State machine states:
    type \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._States\ is (
        \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_0\, 
        \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_1\, 
        \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_2\, 
        \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_3\, 
        \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_4\, 
        \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_5\, 
        \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_6\);
    -- Signals:
    Signal \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._Finished\: boolean := false;
    Signal \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).indexObject.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.0\: boolean := false;
    Signal \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).indexObject.parameter.Out.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.1\: boolean := false;
    Signal \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).indexObject.parameter.Out.2\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.2\: boolean := false;
    Signal \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._Started\: boolean := false;
    Signal \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.input.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Finished.0\: boolean := false;
    Signal \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Finished.1\: boolean := false;
    Signal \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Finished.2\: boolean := false;
    Signal \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).return.0\: boolean := false;
    Signal \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).return.1\: boolean := false;
    Signal \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).return.2\: boolean := false;
    -- System.Void Hast.TestInputs.Various.ParallelCases::WhenAllWhenAnyAwaitedTasks(System.UInt32).0 declarations end


    -- System.Void Hast.TestInputs.Various.ParallelCases::ObjectUsingTasks(System.UInt32).0 declarations start
    -- State machine states:
    type \ParallelCases::ObjectUsingTasks(UInt32).0._States\ is (
        \ParallelCases::ObjectUsingTasks(UInt32).0._State_0\, 
        \ParallelCases::ObjectUsingTasks(UInt32).0._State_1\, 
        \ParallelCases::ObjectUsingTasks(UInt32).0._State_2\, 
        \ParallelCases::ObjectUsingTasks(UInt32).0._State_3\, 
        \ParallelCases::ObjectUsingTasks(UInt32).0._State_4\, 
        \ParallelCases::ObjectUsingTasks(UInt32).0._State_5\);
    -- Signals:
    Signal \ParallelCases::ObjectUsingTasks(UInt32).0._Finished\: boolean := false;
    Signal \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).indexObject.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Started.0\: boolean := false;
    Signal \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).indexObject.parameter.Out.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Started.1\: boolean := false;
    Signal \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).indexObject.parameter.Out.2\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Started.2\: boolean := false;
    Signal \ParallelCases::ObjectUsingTasks(UInt32).0._Started\: boolean := false;
    Signal \ParallelCases::ObjectUsingTasks(UInt32).0.input.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Finished.0\: boolean := false;
    Signal \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Finished.1\: boolean := false;
    Signal \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Finished.2\: boolean := false;
    Signal \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).return.0\: boolean := false;
    Signal \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).return.1\: boolean := false;
    Signal \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).return.2\: boolean := false;
    -- System.Void Hast.TestInputs.Various.ParallelCases::ObjectUsingTasks(System.UInt32).0 declarations end


    -- System.Void Hast.TestInputs.Various.UnaryCases::IncrementDecrement(System.Int32).0 declarations start
    -- State machine states:
    type \UnaryCases::IncrementDecrement(Int32).0._States\ is (
        \UnaryCases::IncrementDecrement(Int32).0._State_0\, 
        \UnaryCases::IncrementDecrement(Int32).0._State_1\, 
        \UnaryCases::IncrementDecrement(Int32).0._State_2\, 
        \UnaryCases::IncrementDecrement(Int32).0._State_3\, 
        \UnaryCases::IncrementDecrement(Int32).0._State_4\);
    -- Signals:
    Signal \UnaryCases::IncrementDecrement(Int32).0._Finished\: boolean := false;
    Signal \UnaryCases::IncrementDecrement(Int32).0._Started\: boolean := false;
    Signal \UnaryCases::IncrementDecrement(Int32).0.input.parameter.In\: signed(31 downto 0) := to_signed(0, 32);
    -- System.Void Hast.TestInputs.Various.UnaryCases::IncrementDecrement(System.Int32).0 declarations end


    -- System.Void Hast::ExternalInvocationProxy() declarations start
    -- Signals:
    Signal \FinishedInternal\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().RootClass::VirtualMethod(Int32)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1()._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Interface1Method2()._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Interface2Method1()._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1()._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2()._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::NonVirtualNonInterfaceMehod()._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().StaticClass::StaticMethod()._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().UnusedDeclarations::UnusedMethod()._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().StaticReference::StaticClassUsingMethod()._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ArrayUsingCases::PassArrayToConstructor()._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ArrayUsingCases::PassArrayFromMethod()._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().CastingCases::NumberCasting(Int16,Int16)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantValuedVariables(Int32)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantPassingToMethod(Int32)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantPassingToObject()._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().LoopCases::BreakInLoop(Int32)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().LoopCases::BreakInLoopInLoop(Int32)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ObjectUsingCases::NullUsage()._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ObjectUsingCases::VoidReturn(Int32)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ParallelCases::ObjectUsingTasks(UInt32)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().UnaryCases::IncrementDecrement(Int32)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().RootClass::VirtualMethod(Int32)._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1()._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Interface1Method2()._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Interface2Method1()._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1()._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2()._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::NonVirtualNonInterfaceMehod()._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().StaticClass::StaticMethod()._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().UnusedDeclarations::UnusedMethod()._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().StaticReference::StaticClassUsingMethod()._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ArrayUsingCases::PassArrayToConstructor()._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ArrayUsingCases::PassArrayFromMethod()._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().CastingCases::NumberCasting(Int16,Int16)._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantValuedVariables(Int32)._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantPassingToMethod(Int32)._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantPassingToObject()._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().LoopCases::BreakInLoop(Int32)._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().LoopCases::BreakInLoopInLoop(Int32)._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ObjectUsingCases::NullUsage()._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ObjectUsingCases::VoidReturn(Int32)._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32)._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().ParallelCases::ObjectUsingTasks(UInt32)._Finished.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().UnaryCases::IncrementDecrement(Int32)._Finished.0\: boolean := false;
    -- System.Void Hast::ExternalInvocationProxy() declarations end


    -- \System.Void Hast::InternalInvocationProxy()._CommonDeclarations\ declarations start
    type \InternalInvocationProxy_boolean_Array\ is array (integer range <>) of boolean;
    type \Hast::InternalInvocationProxy()._RunningStates\ is (
        WaitingForStarted, 
        WaitingForFinished, 
        AfterFinished);
    -- \System.Void Hast::InternalInvocationProxy()._CommonDeclarations\ declarations end

begin 

    -- System.Void Hast.TestInputs.ClassStructure1.RootClass::VirtualMethod(System.Int32).0 state machine start
    \RootClass::VirtualMethod(Int32).0._StateMachine\: process (\Clock\) 
        Variable \RootClass::VirtualMethod(Int32).0._State\: \RootClass::VirtualMethod(Int32).0._States\ := \RootClass::VirtualMethod(Int32).0._State_0\;
        Variable \RootClass::VirtualMethod(Int32).0.input\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \RootClass::VirtualMethod(Int32).0._Finished\ <= false;
                \RootClass::VirtualMethod(Int32).0._State\ := \RootClass::VirtualMethod(Int32).0._State_0\;
                \RootClass::VirtualMethod(Int32).0.input\ := to_signed(0, 32);
            else 
                case \RootClass::VirtualMethod(Int32).0._State\ is 
                    when \RootClass::VirtualMethod(Int32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\RootClass::VirtualMethod(Int32).0._Started\ = true) then 
                            \RootClass::VirtualMethod(Int32).0._State\ := \RootClass::VirtualMethod(Int32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RootClass::VirtualMethod(Int32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\RootClass::VirtualMethod(Int32).0._Started\ = true) then 
                            \RootClass::VirtualMethod(Int32).0._Finished\ <= true;
                        else 
                            \RootClass::VirtualMethod(Int32).0._Finished\ <= false;
                            \RootClass::VirtualMethod(Int32).0._State\ := \RootClass::VirtualMethod(Int32).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \RootClass::VirtualMethod(Int32).0._State_2\ => 
                        \RootClass::VirtualMethod(Int32).0.input\ := \RootClass::VirtualMethod(Int32).0.input.parameter.In\;
                        \RootClass::VirtualMethod(Int32).0._State\ := \RootClass::VirtualMethod(Int32).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.ClassStructure1.RootClass::VirtualMethod(System.Int32).0 state machine end


    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0 state machine start
    \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._StateMachine\: process (\Clock\) 
        Variable \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._State\: \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._States\ := \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._State_0\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._Finished\ <= false;
                \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0.ComplexTypeHierarchy::PrivateMethod()._Started.0\ <= false;
                \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._State\ := \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._State_0\;
            else 
                case \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._State\ is 
                    when \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._Started\ = true) then 
                            \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._State\ := \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._Started\ = true) then 
                            \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._Finished\ <= true;
                        else 
                            \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._Finished\ <= false;
                            \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._State\ := \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._State_2\ => 
                        -- Starting state machine invocation for the following method: System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::PrivateMethod()
                        \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0.ComplexTypeHierarchy::PrivateMethod()._Started.0\ <= true;
                        \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._State\ := \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::PrivateMethod()
                        if (\ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0.ComplexTypeHierarchy::PrivateMethod()._Started.0\ = \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0.ComplexTypeHierarchy::PrivateMethod()._Finished.0\) then 
                            \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0.ComplexTypeHierarchy::PrivateMethod()._Started.0\ <= false;
                            \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._State\ := \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0 state machine end


    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Interface1Method2().0 state machine start
    \ComplexTypeHierarchy::Interface1Method2().0._StateMachine\: process (\Clock\) 
        Variable \ComplexTypeHierarchy::Interface1Method2().0._State\: \ComplexTypeHierarchy::Interface1Method2().0._States\ := \ComplexTypeHierarchy::Interface1Method2().0._State_0\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ComplexTypeHierarchy::Interface1Method2().0._Finished\ <= false;
                \ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::PrivateMethod()._Started.0\ <= false;
                \ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::StaticMethod()._Started.0\ <= false;
                \ComplexTypeHierarchy::Interface1Method2().0._State\ := \ComplexTypeHierarchy::Interface1Method2().0._State_0\;
            else 
                case \ComplexTypeHierarchy::Interface1Method2().0._State\ is 
                    when \ComplexTypeHierarchy::Interface1Method2().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ComplexTypeHierarchy::Interface1Method2().0._Started\ = true) then 
                            \ComplexTypeHierarchy::Interface1Method2().0._State\ := \ComplexTypeHierarchy::Interface1Method2().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ComplexTypeHierarchy::Interface1Method2().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ComplexTypeHierarchy::Interface1Method2().0._Started\ = true) then 
                            \ComplexTypeHierarchy::Interface1Method2().0._Finished\ <= true;
                        else 
                            \ComplexTypeHierarchy::Interface1Method2().0._Finished\ <= false;
                            \ComplexTypeHierarchy::Interface1Method2().0._State\ := \ComplexTypeHierarchy::Interface1Method2().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ComplexTypeHierarchy::Interface1Method2().0._State_2\ => 
                        -- Starting state machine invocation for the following method: System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::PrivateMethod()
                        \ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::PrivateMethod()._Started.0\ <= true;
                        \ComplexTypeHierarchy::Interface1Method2().0._State\ := \ComplexTypeHierarchy::Interface1Method2().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ComplexTypeHierarchy::Interface1Method2().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::PrivateMethod()
                        if (\ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::PrivateMethod()._Started.0\ = \ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::PrivateMethod()._Finished.0\) then 
                            \ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::PrivateMethod()._Started.0\ <= false;
                            -- Starting state machine invocation for the following method: System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::StaticMethod()
                            \ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::StaticMethod()._Started.0\ <= true;
                            \ComplexTypeHierarchy::Interface1Method2().0._State\ := \ComplexTypeHierarchy::Interface1Method2().0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ComplexTypeHierarchy::Interface1Method2().0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::StaticMethod()
                        if (\ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::StaticMethod()._Started.0\ = \ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::StaticMethod()._Finished.0\) then 
                            \ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::StaticMethod()._Started.0\ <= false;
                            \ComplexTypeHierarchy::Interface1Method2().0._State\ := \ComplexTypeHierarchy::Interface1Method2().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Interface1Method2().0 state machine end


    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Interface2Method1().0 state machine start
    \ComplexTypeHierarchy::Interface2Method1().0._StateMachine\: process (\Clock\) 
        Variable \ComplexTypeHierarchy::Interface2Method1().0._State\: \ComplexTypeHierarchy::Interface2Method1().0._States\ := \ComplexTypeHierarchy::Interface2Method1().0._State_0\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ComplexTypeHierarchy::Interface2Method1().0._Finished\ <= false;
                \ComplexTypeHierarchy::Interface2Method1().0.ComplexTypeHierarchy::BaseInterfaceMethod2()._Started.0\ <= false;
                \ComplexTypeHierarchy::Interface2Method1().0._State\ := \ComplexTypeHierarchy::Interface2Method1().0._State_0\;
            else 
                case \ComplexTypeHierarchy::Interface2Method1().0._State\ is 
                    when \ComplexTypeHierarchy::Interface2Method1().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ComplexTypeHierarchy::Interface2Method1().0._Started\ = true) then 
                            \ComplexTypeHierarchy::Interface2Method1().0._State\ := \ComplexTypeHierarchy::Interface2Method1().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ComplexTypeHierarchy::Interface2Method1().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ComplexTypeHierarchy::Interface2Method1().0._Started\ = true) then 
                            \ComplexTypeHierarchy::Interface2Method1().0._Finished\ <= true;
                        else 
                            \ComplexTypeHierarchy::Interface2Method1().0._Finished\ <= false;
                            \ComplexTypeHierarchy::Interface2Method1().0._State\ := \ComplexTypeHierarchy::Interface2Method1().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ComplexTypeHierarchy::Interface2Method1().0._State_2\ => 
                        -- Starting state machine invocation for the following method: System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::BaseInterfaceMethod2()
                        \ComplexTypeHierarchy::Interface2Method1().0.ComplexTypeHierarchy::BaseInterfaceMethod2()._Started.0\ <= true;
                        \ComplexTypeHierarchy::Interface2Method1().0._State\ := \ComplexTypeHierarchy::Interface2Method1().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ComplexTypeHierarchy::Interface2Method1().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::BaseInterfaceMethod2()
                        if (\ComplexTypeHierarchy::Interface2Method1().0.ComplexTypeHierarchy::BaseInterfaceMethod2()._Started.0\ = \ComplexTypeHierarchy::Interface2Method1().0.ComplexTypeHierarchy::BaseInterfaceMethod2()._Finished.0\) then 
                            \ComplexTypeHierarchy::Interface2Method1().0.ComplexTypeHierarchy::BaseInterfaceMethod2()._Started.0\ <= false;
                            \ComplexTypeHierarchy::Interface2Method1().0._State\ := \ComplexTypeHierarchy::Interface2Method1().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Interface2Method1().0 state machine end


    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0 state machine start
    \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._StateMachine\: process (\Clock\) 
        Variable \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._State\: \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._States\ := \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._State_0\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._Finished\ <= false;
                \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._State\ := \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._State_0\;
            else 
                case \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._State\ is 
                    when \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._Started\ = true) then 
                            \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._State\ := \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._Started\ = true) then 
                            \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._Finished\ <= true;
                        else 
                            \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._Finished\ <= false;
                            \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._State\ := \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._State_2\ => 
                        \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._State\ := \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0 state machine end


    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::BaseInterfaceMethod2().0 state machine start
    \ComplexTypeHierarchy::BaseInterfaceMethod2().0._StateMachine\: process (\Clock\) 
        Variable \ComplexTypeHierarchy::BaseInterfaceMethod2().0._State\: \ComplexTypeHierarchy::BaseInterfaceMethod2().0._States\ := \ComplexTypeHierarchy::BaseInterfaceMethod2().0._State_0\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ComplexTypeHierarchy::BaseInterfaceMethod2().0._Finished\ <= false;
                \ComplexTypeHierarchy::BaseInterfaceMethod2().0.ComplexTypeHierarchy::StaticMethod()._Started.0\ <= false;
                \ComplexTypeHierarchy::BaseInterfaceMethod2().0._State\ := \ComplexTypeHierarchy::BaseInterfaceMethod2().0._State_0\;
            else 
                case \ComplexTypeHierarchy::BaseInterfaceMethod2().0._State\ is 
                    when \ComplexTypeHierarchy::BaseInterfaceMethod2().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ComplexTypeHierarchy::BaseInterfaceMethod2().0._Started\ = true) then 
                            \ComplexTypeHierarchy::BaseInterfaceMethod2().0._State\ := \ComplexTypeHierarchy::BaseInterfaceMethod2().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ComplexTypeHierarchy::BaseInterfaceMethod2().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ComplexTypeHierarchy::BaseInterfaceMethod2().0._Started\ = true) then 
                            \ComplexTypeHierarchy::BaseInterfaceMethod2().0._Finished\ <= true;
                        else 
                            \ComplexTypeHierarchy::BaseInterfaceMethod2().0._Finished\ <= false;
                            \ComplexTypeHierarchy::BaseInterfaceMethod2().0._State\ := \ComplexTypeHierarchy::BaseInterfaceMethod2().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ComplexTypeHierarchy::BaseInterfaceMethod2().0._State_2\ => 
                        -- Starting state machine invocation for the following method: System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::StaticMethod()
                        \ComplexTypeHierarchy::BaseInterfaceMethod2().0.ComplexTypeHierarchy::StaticMethod()._Started.0\ <= true;
                        \ComplexTypeHierarchy::BaseInterfaceMethod2().0._State\ := \ComplexTypeHierarchy::BaseInterfaceMethod2().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ComplexTypeHierarchy::BaseInterfaceMethod2().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::StaticMethod()
                        if (\ComplexTypeHierarchy::BaseInterfaceMethod2().0.ComplexTypeHierarchy::StaticMethod()._Started.0\ = \ComplexTypeHierarchy::BaseInterfaceMethod2().0.ComplexTypeHierarchy::StaticMethod()._Finished.0\) then 
                            \ComplexTypeHierarchy::BaseInterfaceMethod2().0.ComplexTypeHierarchy::StaticMethod()._Started.0\ <= false;
                            \ComplexTypeHierarchy::BaseInterfaceMethod2().0._State\ := \ComplexTypeHierarchy::BaseInterfaceMethod2().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::BaseInterfaceMethod2().0 state machine end


    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0 state machine start
    \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._StateMachine\: process (\Clock\) 
        Variable \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._State\: \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._States\ := \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._State_0\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._Finished\ <= false;
                \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0.ComplexTypeHierarchy::PrivateMethod()._Started.0\ <= false;
                \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._State\ := \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._State_0\;
            else 
                case \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._State\ is 
                    when \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._Started\ = true) then 
                            \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._State\ := \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._Started\ = true) then 
                            \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._Finished\ <= true;
                        else 
                            \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._Finished\ <= false;
                            \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._State\ := \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._State_2\ => 
                        -- Starting state machine invocation for the following method: System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::PrivateMethod()
                        \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0.ComplexTypeHierarchy::PrivateMethod()._Started.0\ <= true;
                        \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._State\ := \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::PrivateMethod()
                        if (\ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0.ComplexTypeHierarchy::PrivateMethod()._Started.0\ = \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0.ComplexTypeHierarchy::PrivateMethod()._Finished.0\) then 
                            \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0.ComplexTypeHierarchy::PrivateMethod()._Started.0\ <= false;
                            \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._State\ := \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0 state machine end


    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::PrivateMethod().0 state machine start
    \ComplexTypeHierarchy::PrivateMethod().0._StateMachine\: process (\Clock\) 
        Variable \ComplexTypeHierarchy::PrivateMethod().0._State\: \ComplexTypeHierarchy::PrivateMethod().0._States\ := \ComplexTypeHierarchy::PrivateMethod().0._State_0\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ComplexTypeHierarchy::PrivateMethod().0._Finished\ <= false;
                \ComplexTypeHierarchy::PrivateMethod().0.ComplexTypeHierarchy::StaticMethod()._Started.0\ <= false;
                \ComplexTypeHierarchy::PrivateMethod().0._State\ := \ComplexTypeHierarchy::PrivateMethod().0._State_0\;
            else 
                case \ComplexTypeHierarchy::PrivateMethod().0._State\ is 
                    when \ComplexTypeHierarchy::PrivateMethod().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ComplexTypeHierarchy::PrivateMethod().0._Started\ = true) then 
                            \ComplexTypeHierarchy::PrivateMethod().0._State\ := \ComplexTypeHierarchy::PrivateMethod().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ComplexTypeHierarchy::PrivateMethod().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ComplexTypeHierarchy::PrivateMethod().0._Started\ = true) then 
                            \ComplexTypeHierarchy::PrivateMethod().0._Finished\ <= true;
                        else 
                            \ComplexTypeHierarchy::PrivateMethod().0._Finished\ <= false;
                            \ComplexTypeHierarchy::PrivateMethod().0._State\ := \ComplexTypeHierarchy::PrivateMethod().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ComplexTypeHierarchy::PrivateMethod().0._State_2\ => 
                        -- Starting state machine invocation for the following method: System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::StaticMethod()
                        \ComplexTypeHierarchy::PrivateMethod().0.ComplexTypeHierarchy::StaticMethod()._Started.0\ <= true;
                        \ComplexTypeHierarchy::PrivateMethod().0._State\ := \ComplexTypeHierarchy::PrivateMethod().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ComplexTypeHierarchy::PrivateMethod().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::StaticMethod()
                        if (\ComplexTypeHierarchy::PrivateMethod().0.ComplexTypeHierarchy::StaticMethod()._Started.0\ = \ComplexTypeHierarchy::PrivateMethod().0.ComplexTypeHierarchy::StaticMethod()._Finished.0\) then 
                            \ComplexTypeHierarchy::PrivateMethod().0.ComplexTypeHierarchy::StaticMethod()._Started.0\ <= false;
                            \ComplexTypeHierarchy::PrivateMethod().0._State\ := \ComplexTypeHierarchy::PrivateMethod().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::PrivateMethod().0 state machine end


    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::StaticMethod().0 state machine start
    \ComplexTypeHierarchy::StaticMethod().0._StateMachine\: process (\Clock\) 
        Variable \ComplexTypeHierarchy::StaticMethod().0._State\: \ComplexTypeHierarchy::StaticMethod().0._States\ := \ComplexTypeHierarchy::StaticMethod().0._State_0\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ComplexTypeHierarchy::StaticMethod().0._Finished\ <= false;
                \ComplexTypeHierarchy::StaticMethod().0._State\ := \ComplexTypeHierarchy::StaticMethod().0._State_0\;
            else 
                case \ComplexTypeHierarchy::StaticMethod().0._State\ is 
                    when \ComplexTypeHierarchy::StaticMethod().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ComplexTypeHierarchy::StaticMethod().0._Started\ = true) then 
                            \ComplexTypeHierarchy::StaticMethod().0._State\ := \ComplexTypeHierarchy::StaticMethod().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ComplexTypeHierarchy::StaticMethod().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ComplexTypeHierarchy::StaticMethod().0._Started\ = true) then 
                            \ComplexTypeHierarchy::StaticMethod().0._Finished\ <= true;
                        else 
                            \ComplexTypeHierarchy::StaticMethod().0._Finished\ <= false;
                            \ComplexTypeHierarchy::StaticMethod().0._State\ := \ComplexTypeHierarchy::StaticMethod().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ComplexTypeHierarchy::StaticMethod().0._State_2\ => 
                        \ComplexTypeHierarchy::StaticMethod().0._State\ := \ComplexTypeHierarchy::StaticMethod().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::StaticMethod().0 state machine end


    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.StaticClass::StaticMethod().0 state machine start
    \StaticClass::StaticMethod().0._StateMachine\: process (\Clock\) 
        Variable \StaticClass::StaticMethod().0._State\: \StaticClass::StaticMethod().0._States\ := \StaticClass::StaticMethod().0._State_0\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \StaticClass::StaticMethod().0._Finished\ <= false;
                \StaticClass::StaticMethod().0._State\ := \StaticClass::StaticMethod().0._State_0\;
            else 
                case \StaticClass::StaticMethod().0._State\ is 
                    when \StaticClass::StaticMethod().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\StaticClass::StaticMethod().0._Started\ = true) then 
                            \StaticClass::StaticMethod().0._State\ := \StaticClass::StaticMethod().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \StaticClass::StaticMethod().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\StaticClass::StaticMethod().0._Started\ = true) then 
                            \StaticClass::StaticMethod().0._Finished\ <= true;
                        else 
                            \StaticClass::StaticMethod().0._Finished\ <= false;
                            \StaticClass::StaticMethod().0._State\ := \StaticClass::StaticMethod().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \StaticClass::StaticMethod().0._State_2\ => 
                        \StaticClass::StaticMethod().0._State\ := \StaticClass::StaticMethod().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.StaticClass::StaticMethod().0 state machine end


    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.UnusedDeclarations::UnusedMethod().0 state machine start
    \UnusedDeclarations::UnusedMethod().0._StateMachine\: process (\Clock\) 
        Variable \UnusedDeclarations::UnusedMethod().0._State\: \UnusedDeclarations::UnusedMethod().0._States\ := \UnusedDeclarations::UnusedMethod().0._State_0\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \UnusedDeclarations::UnusedMethod().0._Finished\ <= false;
                \UnusedDeclarations::UnusedMethod().0._State\ := \UnusedDeclarations::UnusedMethod().0._State_0\;
            else 
                case \UnusedDeclarations::UnusedMethod().0._State\ is 
                    when \UnusedDeclarations::UnusedMethod().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\UnusedDeclarations::UnusedMethod().0._Started\ = true) then 
                            \UnusedDeclarations::UnusedMethod().0._State\ := \UnusedDeclarations::UnusedMethod().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnusedDeclarations::UnusedMethod().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\UnusedDeclarations::UnusedMethod().0._Started\ = true) then 
                            \UnusedDeclarations::UnusedMethod().0._Finished\ <= true;
                        else 
                            \UnusedDeclarations::UnusedMethod().0._Finished\ <= false;
                            \UnusedDeclarations::UnusedMethod().0._State\ := \UnusedDeclarations::UnusedMethod().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnusedDeclarations::UnusedMethod().0._State_2\ => 
                        \UnusedDeclarations::UnusedMethod().0._State\ := \UnusedDeclarations::UnusedMethod().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.UnusedDeclarations::UnusedMethod().0 state machine end


    -- System.Void Hast.TestInputs.ClassStructure2.StaticReference::StaticClassUsingMethod().0 state machine start
    \StaticReference::StaticClassUsingMethod().0._StateMachine\: process (\Clock\) 
        Variable \StaticReference::StaticClassUsingMethod().0._State\: \StaticReference::StaticClassUsingMethod().0._States\ := \StaticReference::StaticClassUsingMethod().0._State_0\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \StaticReference::StaticClassUsingMethod().0._Finished\ <= false;
                \StaticReference::StaticClassUsingMethod().0.StaticClass::StaticMethod()._Started.0\ <= false;
                \StaticReference::StaticClassUsingMethod().0._State\ := \StaticReference::StaticClassUsingMethod().0._State_0\;
            else 
                case \StaticReference::StaticClassUsingMethod().0._State\ is 
                    when \StaticReference::StaticClassUsingMethod().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\StaticReference::StaticClassUsingMethod().0._Started\ = true) then 
                            \StaticReference::StaticClassUsingMethod().0._State\ := \StaticReference::StaticClassUsingMethod().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \StaticReference::StaticClassUsingMethod().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\StaticReference::StaticClassUsingMethod().0._Started\ = true) then 
                            \StaticReference::StaticClassUsingMethod().0._Finished\ <= true;
                        else 
                            \StaticReference::StaticClassUsingMethod().0._Finished\ <= false;
                            \StaticReference::StaticClassUsingMethod().0._State\ := \StaticReference::StaticClassUsingMethod().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \StaticReference::StaticClassUsingMethod().0._State_2\ => 
                        -- Starting state machine invocation for the following method: System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.StaticClass::StaticMethod()
                        \StaticReference::StaticClassUsingMethod().0.StaticClass::StaticMethod()._Started.0\ <= true;
                        \StaticReference::StaticClassUsingMethod().0._State\ := \StaticReference::StaticClassUsingMethod().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \StaticReference::StaticClassUsingMethod().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.StaticClass::StaticMethod()
                        if (\StaticReference::StaticClassUsingMethod().0.StaticClass::StaticMethod()._Started.0\ = \StaticReference::StaticClassUsingMethod().0.StaticClass::StaticMethod()._Finished.0\) then 
                            \StaticReference::StaticClassUsingMethod().0.StaticClass::StaticMethod()._Started.0\ <= false;
                            \StaticReference::StaticClassUsingMethod().0._State\ := \StaticReference::StaticClassUsingMethod().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.ClassStructure2.StaticReference::StaticClassUsingMethod().0 state machine end


    -- System.Void Hast.TestInputs.Various.ArrayUsingCases/ArrayHolder::.ctor(System.Int32[]).0 state machine start
    \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._StateMachine\: process (\Clock\) 
        Variable \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._State\: \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._States\ := \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._State_0\;
        Variable \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0.this\: \Hast.TestInputs.Various.ArrayUsingCases/ArrayHolder\;
        Variable \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0.array\: \signed32_Array\(0 to 4) := (others => to_signed(0, 32));
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._Finished\ <= false;
                \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0.array.parameter.Out\ <= (others => to_signed(0, 32));
                \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._State\ := \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._State_0\;
                \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0.array\ := (others => to_signed(0, 32));
            else 
                case \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._State\ is 
                    when \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._Started\ = true) then 
                            \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._State\ := \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._Started\ = true) then 
                            \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._Finished\ <= true;
                        else 
                            \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._Finished\ <= false;
                            \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._State\ := \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0.this.parameter.Out\ <= \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0.this\;
                        \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0.array.parameter.Out\ <= \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0.array\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._State_2\ => 
                        \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0.this\ := \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0.this.parameter.In\;
                        \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0.array\ := \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0.array.parameter.In\;
                        \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0.this\.\Array\ := \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0.array\;
                        \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._State\ := \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.Various.ArrayUsingCases/ArrayHolder::.ctor(System.Int32[]).0 state machine end


    -- System.Void Hast.TestInputs.Various.ArrayUsingCases::PassArrayToConstructor().0 state machine start
    \ArrayUsingCases::PassArrayToConstructor().0._StateMachine\: process (\Clock\) 
        Variable \ArrayUsingCases::PassArrayToConstructor().0._State\: \ArrayUsingCases::PassArrayToConstructor().0._States\ := \ArrayUsingCases::PassArrayToConstructor().0._State_0\;
        Variable \ArrayUsingCases::PassArrayToConstructor().0.array\: \signed32_Array\(0 to 4) := (others => to_signed(0, 32));
        Variable \ArrayUsingCases::PassArrayToConstructor().0.arrayHolder\: \Hast.TestInputs.Various.ArrayUsingCases/ArrayHolder\;
        Variable \ArrayUsingCases::PassArrayToConstructor().0.num\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ArrayUsingCases::PassArrayToConstructor().0._Finished\ <= false;
                \ArrayUsingCases::PassArrayToConstructor().0.ArrayUsingCases/ArrayHolder::.ctor(Int32[]).array.parameter.Out.0\ <= (others => to_signed(0, 32));
                \ArrayUsingCases::PassArrayToConstructor().0.ArrayUsingCases/ArrayHolder::.ctor(Int32[])._Started.0\ <= false;
                \ArrayUsingCases::PassArrayToConstructor().0._State\ := \ArrayUsingCases::PassArrayToConstructor().0._State_0\;
                \ArrayUsingCases::PassArrayToConstructor().0.array\ := (others => to_signed(0, 32));
                \ArrayUsingCases::PassArrayToConstructor().0.num\ := to_signed(0, 32);
            else 
                case \ArrayUsingCases::PassArrayToConstructor().0._State\ is 
                    when \ArrayUsingCases::PassArrayToConstructor().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ArrayUsingCases::PassArrayToConstructor().0._Started\ = true) then 
                            \ArrayUsingCases::PassArrayToConstructor().0._State\ := \ArrayUsingCases::PassArrayToConstructor().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ArrayUsingCases::PassArrayToConstructor().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ArrayUsingCases::PassArrayToConstructor().0._Started\ = true) then 
                            \ArrayUsingCases::PassArrayToConstructor().0._Finished\ <= true;
                        else 
                            \ArrayUsingCases::PassArrayToConstructor().0._Finished\ <= false;
                            \ArrayUsingCases::PassArrayToConstructor().0._State\ := \ArrayUsingCases::PassArrayToConstructor().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ArrayUsingCases::PassArrayToConstructor().0._State_2\ => 
                        \ArrayUsingCases::PassArrayToConstructor().0.array\ := (others => to_signed(0, 32));
                        -- Initializing record fields to their defaults.
                        \ArrayUsingCases::PassArrayToConstructor().0.arrayHolder\.\IsNull\ := false;
                        \ArrayUsingCases::PassArrayToConstructor().0.arrayHolder\.\Array\ := (others => to_signed(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Hast.TestInputs.Various.ArrayUsingCases/ArrayHolder::.ctor(System.Int32[])
                        \ArrayUsingCases::PassArrayToConstructor().0.ArrayUsingCases/ArrayHolder::.ctor(Int32[]).this.parameter.Out.0\ <= \ArrayUsingCases::PassArrayToConstructor().0.arrayHolder\;
                        \ArrayUsingCases::PassArrayToConstructor().0.ArrayUsingCases/ArrayHolder::.ctor(Int32[]).array.parameter.Out.0\ <= \ArrayUsingCases::PassArrayToConstructor().0.array\;
                        \ArrayUsingCases::PassArrayToConstructor().0.ArrayUsingCases/ArrayHolder::.ctor(Int32[])._Started.0\ <= true;
                        \ArrayUsingCases::PassArrayToConstructor().0._State\ := \ArrayUsingCases::PassArrayToConstructor().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ArrayUsingCases::PassArrayToConstructor().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.TestInputs.Various.ArrayUsingCases/ArrayHolder::.ctor(System.Int32[])
                        if (\ArrayUsingCases::PassArrayToConstructor().0.ArrayUsingCases/ArrayHolder::.ctor(Int32[])._Started.0\ = \ArrayUsingCases::PassArrayToConstructor().0.ArrayUsingCases/ArrayHolder::.ctor(Int32[])._Finished.0\) then 
                            \ArrayUsingCases::PassArrayToConstructor().0.ArrayUsingCases/ArrayHolder::.ctor(Int32[])._Started.0\ <= false;
                            \ArrayUsingCases::PassArrayToConstructor().0.arrayHolder\ := \ArrayUsingCases::PassArrayToConstructor().0.ArrayUsingCases/ArrayHolder::.ctor(Int32[]).this.parameter.In.0\;
                            \ArrayUsingCases::PassArrayToConstructor().0.array\ := \ArrayUsingCases::PassArrayToConstructor().0.ArrayUsingCases/ArrayHolder::.ctor(Int32[]).array.parameter.In.0\;
                            \ArrayUsingCases::PassArrayToConstructor().0.num\ := to_signed(5, 32);
                            \ArrayUsingCases::PassArrayToConstructor().0._State\ := \ArrayUsingCases::PassArrayToConstructor().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.Various.ArrayUsingCases::PassArrayToConstructor().0 state machine end


    -- System.Void Hast.TestInputs.Various.ArrayUsingCases::PassArrayFromMethod().0 state machine start
    \ArrayUsingCases::PassArrayFromMethod().0._StateMachine\: process (\Clock\) 
        Variable \ArrayUsingCases::PassArrayFromMethod().0._State\: \ArrayUsingCases::PassArrayFromMethod().0._States\ := \ArrayUsingCases::PassArrayFromMethod().0._State_0\;
        Variable \ArrayUsingCases::PassArrayFromMethod().0.array\: \signed32_Array\(0 to 4) := (others => to_signed(0, 32));
        Variable \ArrayUsingCases::PassArrayFromMethod().0.return.0\: \signed32_Array\(0 to 4) := (others => to_signed(0, 32));
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ArrayUsingCases::PassArrayFromMethod().0._Finished\ <= false;
                \ArrayUsingCases::PassArrayFromMethod().0.ArrayUsingCases::ArrayProducingMethod(Int32).arrayLength.parameter.Out.0\ <= to_signed(0, 32);
                \ArrayUsingCases::PassArrayFromMethod().0.ArrayUsingCases::ArrayProducingMethod(Int32)._Started.0\ <= false;
                \ArrayUsingCases::PassArrayFromMethod().0._State\ := \ArrayUsingCases::PassArrayFromMethod().0._State_0\;
                \ArrayUsingCases::PassArrayFromMethod().0.array\ := (others => to_signed(0, 32));
                \ArrayUsingCases::PassArrayFromMethod().0.return.0\ := (others => to_signed(0, 32));
            else 
                case \ArrayUsingCases::PassArrayFromMethod().0._State\ is 
                    when \ArrayUsingCases::PassArrayFromMethod().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ArrayUsingCases::PassArrayFromMethod().0._Started\ = true) then 
                            \ArrayUsingCases::PassArrayFromMethod().0._State\ := \ArrayUsingCases::PassArrayFromMethod().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ArrayUsingCases::PassArrayFromMethod().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ArrayUsingCases::PassArrayFromMethod().0._Started\ = true) then 
                            \ArrayUsingCases::PassArrayFromMethod().0._Finished\ <= true;
                        else 
                            \ArrayUsingCases::PassArrayFromMethod().0._Finished\ <= false;
                            \ArrayUsingCases::PassArrayFromMethod().0._State\ := \ArrayUsingCases::PassArrayFromMethod().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ArrayUsingCases::PassArrayFromMethod().0._State_2\ => 
                        -- Starting state machine invocation for the following method: System.Int32[] Hast.TestInputs.Various.ArrayUsingCases::ArrayProducingMethod(System.Int32)
                        \ArrayUsingCases::PassArrayFromMethod().0.ArrayUsingCases::ArrayProducingMethod(Int32).arrayLength.parameter.Out.0\ <= to_signed(5, 32);
                        \ArrayUsingCases::PassArrayFromMethod().0.ArrayUsingCases::ArrayProducingMethod(Int32)._Started.0\ <= true;
                        \ArrayUsingCases::PassArrayFromMethod().0._State\ := \ArrayUsingCases::PassArrayFromMethod().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ArrayUsingCases::PassArrayFromMethod().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Int32[] Hast.TestInputs.Various.ArrayUsingCases::ArrayProducingMethod(System.Int32)
                        if (\ArrayUsingCases::PassArrayFromMethod().0.ArrayUsingCases::ArrayProducingMethod(Int32)._Started.0\ = \ArrayUsingCases::PassArrayFromMethod().0.ArrayUsingCases::ArrayProducingMethod(Int32)._Finished.0\) then 
                            \ArrayUsingCases::PassArrayFromMethod().0.ArrayUsingCases::ArrayProducingMethod(Int32)._Started.0\ <= false;
                            \ArrayUsingCases::PassArrayFromMethod().0.return.0\ := \ArrayUsingCases::PassArrayFromMethod().0.ArrayUsingCases::ArrayProducingMethod(Int32).return.0\;
                            \ArrayUsingCases::PassArrayFromMethod().0.array\ := \ArrayUsingCases::PassArrayFromMethod().0.return.0\;
                            \ArrayUsingCases::PassArrayFromMethod().0._State\ := \ArrayUsingCases::PassArrayFromMethod().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.Various.ArrayUsingCases::PassArrayFromMethod().0 state machine end


    -- System.Int32[] Hast.TestInputs.Various.ArrayUsingCases::ArrayProducingMethod(System.Int32).0 state machine start
    \ArrayUsingCases::ArrayProducingMethod(Int32).0._StateMachine\: process (\Clock\) 
        Variable \ArrayUsingCases::ArrayProducingMethod(Int32).0._State\: \ArrayUsingCases::ArrayProducingMethod(Int32).0._States\ := \ArrayUsingCases::ArrayProducingMethod(Int32).0._State_0\;
        Variable \ArrayUsingCases::ArrayProducingMethod(Int32).0.arrayLength\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ArrayUsingCases::ArrayProducingMethod(Int32).0.array\: \signed32_Array\(0 to 4) := (others => to_signed(0, 32));
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ArrayUsingCases::ArrayProducingMethod(Int32).0._Finished\ <= false;
                \ArrayUsingCases::ArrayProducingMethod(Int32).0.return\ <= (others => to_signed(0, 32));
                \ArrayUsingCases::ArrayProducingMethod(Int32).0._State\ := \ArrayUsingCases::ArrayProducingMethod(Int32).0._State_0\;
                \ArrayUsingCases::ArrayProducingMethod(Int32).0.arrayLength\ := to_signed(0, 32);
                \ArrayUsingCases::ArrayProducingMethod(Int32).0.array\ := (others => to_signed(0, 32));
            else 
                case \ArrayUsingCases::ArrayProducingMethod(Int32).0._State\ is 
                    when \ArrayUsingCases::ArrayProducingMethod(Int32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ArrayUsingCases::ArrayProducingMethod(Int32).0._Started\ = true) then 
                            \ArrayUsingCases::ArrayProducingMethod(Int32).0._State\ := \ArrayUsingCases::ArrayProducingMethod(Int32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ArrayUsingCases::ArrayProducingMethod(Int32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ArrayUsingCases::ArrayProducingMethod(Int32).0._Started\ = true) then 
                            \ArrayUsingCases::ArrayProducingMethod(Int32).0._Finished\ <= true;
                        else 
                            \ArrayUsingCases::ArrayProducingMethod(Int32).0._Finished\ <= false;
                            \ArrayUsingCases::ArrayProducingMethod(Int32).0._State\ := \ArrayUsingCases::ArrayProducingMethod(Int32).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ArrayUsingCases::ArrayProducingMethod(Int32).0._State_2\ => 
                        \ArrayUsingCases::ArrayProducingMethod(Int32).0.arrayLength\ := \ArrayUsingCases::ArrayProducingMethod(Int32).0.arrayLength.parameter.In\;
                        \ArrayUsingCases::ArrayProducingMethod(Int32).0.array\ := (others => to_signed(0, 32));
                        \ArrayUsingCases::ArrayProducingMethod(Int32).0.array\(to_integer(to_signed(3, 32))) := to_signed(10, 32);
                        \ArrayUsingCases::ArrayProducingMethod(Int32).0.return\ <= \ArrayUsingCases::ArrayProducingMethod(Int32).0.array\;
                        \ArrayUsingCases::ArrayProducingMethod(Int32).0._State\ := \ArrayUsingCases::ArrayProducingMethod(Int32).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Int32[] Hast.TestInputs.Various.ArrayUsingCases::ArrayProducingMethod(System.Int32).0 state machine end


    -- System.Void Hast.TestInputs.Various.CastingCases::NumberCasting(System.Int16,System.Int16).0 state machine start
    \CastingCases::NumberCasting(Int16,Int16).0._StateMachine\: process (\Clock\) 
        Variable \CastingCases::NumberCasting(Int16,Int16).0._State\: \CastingCases::NumberCasting(Int16,Int16).0._States\ := \CastingCases::NumberCasting(Int16,Int16).0._State_0\;
        Variable \CastingCases::NumberCasting(Int16,Int16).0.a\: signed(15 downto 0) := to_signed(0, 16);
        Variable \CastingCases::NumberCasting(Int16,Int16).0.b\: signed(15 downto 0) := to_signed(0, 16);
        Variable \CastingCases::NumberCasting(Int16,Int16).0.num\: signed(15 downto 0) := to_signed(0, 16);
        Variable \CastingCases::NumberCasting(Int16,Int16).0.num2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \CastingCases::NumberCasting(Int16,Int16).0.binaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \CastingCases::NumberCasting(Int16,Int16).0.binaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \CastingCases::NumberCasting(Int16,Int16).0._Finished\ <= false;
                \CastingCases::NumberCasting(Int16,Int16).0._State\ := \CastingCases::NumberCasting(Int16,Int16).0._State_0\;
                \CastingCases::NumberCasting(Int16,Int16).0.a\ := to_signed(0, 16);
                \CastingCases::NumberCasting(Int16,Int16).0.b\ := to_signed(0, 16);
                \CastingCases::NumberCasting(Int16,Int16).0.num\ := to_signed(0, 16);
                \CastingCases::NumberCasting(Int16,Int16).0.num2\ := to_signed(0, 32);
                \CastingCases::NumberCasting(Int16,Int16).0.binaryOperationResult.0\ := to_signed(0, 32);
                \CastingCases::NumberCasting(Int16,Int16).0.binaryOperationResult.1\ := to_signed(0, 32);
            else 
                case \CastingCases::NumberCasting(Int16,Int16).0._State\ is 
                    when \CastingCases::NumberCasting(Int16,Int16).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\CastingCases::NumberCasting(Int16,Int16).0._Started\ = true) then 
                            \CastingCases::NumberCasting(Int16,Int16).0._State\ := \CastingCases::NumberCasting(Int16,Int16).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \CastingCases::NumberCasting(Int16,Int16).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\CastingCases::NumberCasting(Int16,Int16).0._Started\ = true) then 
                            \CastingCases::NumberCasting(Int16,Int16).0._Finished\ <= true;
                        else 
                            \CastingCases::NumberCasting(Int16,Int16).0._Finished\ <= false;
                            \CastingCases::NumberCasting(Int16,Int16).0._State\ := \CastingCases::NumberCasting(Int16,Int16).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \CastingCases::NumberCasting(Int16,Int16).0._State_2\ => 
                        \CastingCases::NumberCasting(Int16,Int16).0.a\ := \CastingCases::NumberCasting(Int16,Int16).0.a.parameter.In\;
                        \CastingCases::NumberCasting(Int16,Int16).0.b\ := \CastingCases::NumberCasting(Int16,Int16).0.b.parameter.In\;
                        \CastingCases::NumberCasting(Int16,Int16).0.binaryOperationResult.0\ := signed(resize(\CastingCases::NumberCasting(Int16,Int16).0.a\ * \CastingCases::NumberCasting(Int16,Int16).0.b\, 32));
                        \CastingCases::NumberCasting(Int16,Int16).0.num\ := \CastingCases::NumberCasting(Int16,Int16).0.binaryOperationResult.0\;
                        \CastingCases::NumberCasting(Int16,Int16).0.binaryOperationResult.1\ := resize(\CastingCases::NumberCasting(Int16,Int16).0.a\ * \CastingCases::NumberCasting(Int16,Int16).0.b\, 32);
                        \CastingCases::NumberCasting(Int16,Int16).0.num2\ := (\CastingCases::NumberCasting(Int16,Int16).0.binaryOperationResult.1\);
                        \CastingCases::NumberCasting(Int16,Int16).0._State\ := \CastingCases::NumberCasting(Int16,Int16).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.Various.CastingCases::NumberCasting(System.Int16,System.Int16).0 state machine end


    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32[]).0 state machine start
    \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._StateMachine\: process (\Clock\) 
        Variable \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._State\: \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._States\ := \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._State_0\;
        Variable \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.this\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
        Variable \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.array\: \unsigned32_Array\(0 to 4) := (others => to_unsigned(0, 32));
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._Finished\ <= false;
                \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.array.parameter.Out\ <= (others => to_unsigned(0, 32));
                \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._State\ := \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._State_0\;
                \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.array\ := (others => to_unsigned(0, 32));
            else 
                case \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._State\ is 
                    when \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._Started\ = true) then 
                            \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._State\ := \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._Started\ = true) then 
                            \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._Finished\ <= true;
                        else 
                            \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._Finished\ <= false;
                            \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._State\ := \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.this.parameter.Out\ <= \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.this\;
                        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.array.parameter.Out\ <= \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.array\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._State_2\ => 
                        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.this\ := \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.this.parameter.In\;
                        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.array\ := \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.array.parameter.In\;
                        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.this\.\ArrayLength\ := to_unsigned(5, 32);
                        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.this\.\ArrayLengthCopy\ := to_unsigned(160, 32);
                        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.this\.\NonSubstitutableArrayLengthCopy\ := to_unsigned(160, 32);
                        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.this\.\Array\ := (others => to_unsigned(0, 32));
                        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._State\ := \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32[]).0 state machine end


    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32).0 state machine start
    \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._StateMachine\: process (\Clock\) 
        Variable \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._State\: \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._States\ := \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._State_0\;
        Variable \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0.this\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
        Variable \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0.size\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0.conditional109a0d002e7b6a56b1572efc4bfd5a39a757d5e88ee9e1fdaf585033fba598d2\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._Finished\ <= false;
                \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._State\ := \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._State_0\;
                \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0.size\ := to_unsigned(0, 32);
                \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0.conditional109a0d002e7b6a56b1572efc4bfd5a39a757d5e88ee9e1fdaf585033fba598d2\ := to_unsigned(0, 32);
            else 
                case \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._State\ is 
                    when \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._Started\ = true) then 
                            \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._State\ := \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._Started\ = true) then 
                            \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._Finished\ <= true;
                        else 
                            \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._Finished\ <= false;
                            \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._State\ := \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0.this.parameter.Out\ <= \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0.this\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._State_2\ => 
                        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0.this\ := \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0.this.parameter.In\;
                        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0.size\ := \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0.size.parameter.In\;
                        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0.conditional109a0d002e7b6a56b1572efc4bfd5a39a757d5e88ee9e1fdaf585033fba598d2\ := to_unsigned(5, 32);
                        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0.this\.\ArrayLength\ := to_unsigned(5, 32);
                        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0.this\.\ArrayLengthCopy\ := to_unsigned(160, 32);
                        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0.this\.\NonSubstitutableArrayLengthCopy\ := to_unsigned(160, 32);
                        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0.this\.\Array\ := (others => to_unsigned(0, 32));
                        \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._State\ := \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32).0 state machine end


    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1).0 state machine start
    \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._StateMachine\: process (\Clock\) 
        Variable \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._State\: \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._States\ := \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._State_0\;
        Variable \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.this\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
        Variable \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.previous\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._Finished\ <= false;
                \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).array.parameter.Out.0\ <= (others => to_unsigned(0, 32));
                \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Started.0\ <= false;
                \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._State\ := \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._State_0\;
            else 
                case \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._State\ is 
                    when \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._Started\ = true) then 
                            \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._State\ := \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._Started\ = true) then 
                            \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._Finished\ <= true;
                        else 
                            \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._Finished\ <= false;
                            \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._State\ := \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.this.parameter.Out\ <= \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.this\;
                        \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.previous.parameter.Out\ <= \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.previous\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._State_2\ => 
                        \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.this\ := \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.this.parameter.In\;
                        \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.previous\ := \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.previous.parameter.In\;
                        -- Starting state machine invocation for the following method: System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32[])
                        \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).this.parameter.Out.0\ <= \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.this\;
                        \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).array.parameter.Out.0\ <= \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.previous\.\Array\;
                        \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Started.0\ <= true;
                        \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._State\ := \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32[])
                        if (\ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Started.0\ = \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Finished.0\) then 
                            \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Started.0\ <= false;
                            \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.this\ := \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).this.parameter.In.0\;
                            \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.previous\.\Array\ := \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).array.parameter.In.0\;
                            \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._State\ := \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1).0 state machine end


    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder2::.ctor(System.UInt32).0 state machine start
    \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._StateMachine\: process (\Clock\) 
        Variable \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State\: \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._States\ := \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_0\;
        Variable \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.this\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder2\;
        Variable \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.size\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.conditional109a0d002e7b6a56b1572efc4bfd5a39a757d5e88ee9e1fdaf585033fba598d2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.binaryOperationResult.1\: boolean := false;
        Variable \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.binaryOperationResult.2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._Finished\ <= false;
                \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State\ := \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_0\;
                \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.size\ := to_unsigned(0, 32);
                \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.conditional109a0d002e7b6a56b1572efc4bfd5a39a757d5e88ee9e1fdaf585033fba598d2\ := to_unsigned(0, 32);
                \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.binaryOperationResult.0\ := to_unsigned(0, 32);
                \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.binaryOperationResult.1\ := false;
                \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.binaryOperationResult.2\ := to_unsigned(0, 32);
                \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.binaryOperationResult.3\ := to_unsigned(0, 32);
            else 
                case \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State\ is 
                    when \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._Started\ = true) then 
                            \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State\ := \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._Started\ = true) then 
                            \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._Finished\ <= true;
                        else 
                            \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._Finished\ <= false;
                            \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State\ := \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.this.parameter.Out\ <= \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.this\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_2\ => 
                        \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.this\ := \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.this.parameter.In\;
                        \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.size\ := \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.size.parameter.In\;
                        \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State\ := \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_3\ => 
                        -- Waiting for the result to appear in \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.binaryOperationResult.0\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State\ := \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_4\;
                            \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ := \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.binaryOperationResult.0\ := \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.size\ mod to_unsigned(32, 32);
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_4\ => 
                        \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.binaryOperationResult.1\ := \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.binaryOperationResult.0\ = to_unsigned(0, 32);

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_6\ and ends in state \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_6\.
                        --     * The false branch starts in state \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_7\ and ends in state \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_7\.
                        --     * Execution after either branch will continue in the following state: \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_5\.

                        if (\ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.binaryOperationResult.1\) then 
                            \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State\ := \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_6\;
                        else 
                            \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State\ := \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_5\ => 
                        -- State after the if-else which was started in state \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_4\.
                        \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.binaryOperationResult.2\ := shift_right(\ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.size\, to_integer(to_signed(5, 32)));
                        \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.binaryOperationResult.3\ := \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.binaryOperationResult.2\ + \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.conditional109a0d002e7b6a56b1572efc4bfd5a39a757d5e88ee9e1fdaf585033fba598d2\;
                        \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.this\.\ArrayLength\ := \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.binaryOperationResult.3\;
                        \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State\ := \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_6\ => 
                        -- True branch of the if-else started in state \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_4\.
                        \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.conditional109a0d002e7b6a56b1572efc4bfd5a39a757d5e88ee9e1fdaf585033fba598d2\ := to_unsigned(0, 32);
                        -- Going to the state after the if-else which was started in state \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_4\.
                        if (\ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State\ = \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_6\) then 
                            \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State\ := \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_7\ => 
                        -- False branch of the if-else started in state \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_4\.
                        \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.conditional109a0d002e7b6a56b1572efc4bfd5a39a757d5e88ee9e1fdaf585033fba598d2\ := to_unsigned(5, 32);
                        -- Going to the state after the if-else which was started in state \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_4\.
                        if (\ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State\ = \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_7\) then 
                            \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State\ := \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder2::.ctor(System.UInt32).0 state machine end


    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases::ConstantValuedVariables(System.Int32).0 state machine start
    \ConstantsUsingCases::ConstantValuedVariables(Int32).0._StateMachine\: process (\Clock\) 
        Variable \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State\: \ConstantsUsingCases::ConstantValuedVariables(Int32).0._States\ := \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_0\;
        Variable \ConstantsUsingCases::ConstantValuedVariables(Int32).0.input\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ConstantsUsingCases::ConstantValuedVariables(Int32).0.num\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ConstantsUsingCases::ConstantValuedVariables(Int32).0.num2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ConstantsUsingCases::ConstantValuedVariables(Int32).0.num3\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ConstantsUsingCases::ConstantValuedVariables(Int32).0.num4\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ConstantsUsingCases::ConstantValuedVariables(Int32).0.array\: \signed32_Array\(0 to 36) := (others => to_signed(0, 32));
        Variable \ConstantsUsingCases::ConstantValuedVariables(Int32).0.num5\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ConstantsUsingCases::ConstantValuedVariables(Int32).0.flag\: boolean := false;
        Variable \ConstantsUsingCases::ConstantValuedVariables(Int32).0.num6\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ConstantsUsingCases::ConstantValuedVariables(Int32).0.flag2\: boolean := false;
        Variable \ConstantsUsingCases::ConstantValuedVariables(Int32).0.binaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ConstantsUsingCases::ConstantValuedVariables(Int32).0.binaryOperationResult.1\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ConstantsUsingCases::ConstantValuedVariables(Int32).0._Finished\ <= false;
                \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State\ := \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_0\;
                \ConstantsUsingCases::ConstantValuedVariables(Int32).0.input\ := to_signed(0, 32);
                \ConstantsUsingCases::ConstantValuedVariables(Int32).0.num\ := to_signed(0, 32);
                \ConstantsUsingCases::ConstantValuedVariables(Int32).0.num2\ := to_signed(0, 32);
                \ConstantsUsingCases::ConstantValuedVariables(Int32).0.num3\ := to_signed(0, 32);
                \ConstantsUsingCases::ConstantValuedVariables(Int32).0.num4\ := to_signed(0, 32);
                \ConstantsUsingCases::ConstantValuedVariables(Int32).0.array\ := (others => to_signed(0, 32));
                \ConstantsUsingCases::ConstantValuedVariables(Int32).0.num5\ := to_signed(0, 32);
                \ConstantsUsingCases::ConstantValuedVariables(Int32).0.flag\ := false;
                \ConstantsUsingCases::ConstantValuedVariables(Int32).0.num6\ := to_signed(0, 32);
                \ConstantsUsingCases::ConstantValuedVariables(Int32).0.flag2\ := false;
                \ConstantsUsingCases::ConstantValuedVariables(Int32).0.binaryOperationResult.0\ := to_signed(0, 32);
                \ConstantsUsingCases::ConstantValuedVariables(Int32).0.binaryOperationResult.1\ := false;
            else 
                case \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State\ is 
                    when \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ConstantsUsingCases::ConstantValuedVariables(Int32).0._Started\ = true) then 
                            \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State\ := \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ConstantsUsingCases::ConstantValuedVariables(Int32).0._Started\ = true) then 
                            \ConstantsUsingCases::ConstantValuedVariables(Int32).0._Finished\ <= true;
                        else 
                            \ConstantsUsingCases::ConstantValuedVariables(Int32).0._Finished\ <= false;
                            \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State\ := \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_2\ => 
                        \ConstantsUsingCases::ConstantValuedVariables(Int32).0.input\ := \ConstantsUsingCases::ConstantValuedVariables(Int32).0.input.parameter.In\;
                        \ConstantsUsingCases::ConstantValuedVariables(Int32).0.num\ := to_signed(4, 32);
                        \ConstantsUsingCases::ConstantValuedVariables(Int32).0.num2\ := to_signed(36, 32);
                        \ConstantsUsingCases::ConstantValuedVariables(Int32).0.num2\ := to_signed(37, 32);
                        \ConstantsUsingCases::ConstantValuedVariables(Int32).0.num3\ := to_signed(148, 32);
                        \ConstantsUsingCases::ConstantValuedVariables(Int32).0.binaryOperationResult.0\ := to_signed(148, 32) + \ConstantsUsingCases::ConstantValuedVariables(Int32).0.input\;
                        \ConstantsUsingCases::ConstantValuedVariables(Int32).0.num4\ := \ConstantsUsingCases::ConstantValuedVariables(Int32).0.binaryOperationResult.0\;
                        \ConstantsUsingCases::ConstantValuedVariables(Int32).0.array\ := (others => to_signed(0, 32));
                        \ConstantsUsingCases::ConstantValuedVariables(Int32).0.num5\ := to_signed(5, 32);
                        \ConstantsUsingCases::ConstantValuedVariables(Int32).0.binaryOperationResult.1\ := \ConstantsUsingCases::ConstantValuedVariables(Int32).0.input\ < to_signed(5, 32);
                        \ConstantsUsingCases::ConstantValuedVariables(Int32).0.flag\ := \ConstantsUsingCases::ConstantValuedVariables(Int32).0.binaryOperationResult.1\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_4\ and ends in state \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_4\.
                        --     * Execution after either branch will continue in the following state: \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_3\.

                        if (\ConstantsUsingCases::ConstantValuedVariables(Int32).0.flag\) then 
                            \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State\ := \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_4\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State\ := \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_3\ => 
                        -- State after the if-else which was started in state \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_2\.
                        \ConstantsUsingCases::ConstantValuedVariables(Int32).0.num6\ := to_signed(153, 32);
                        \ConstantsUsingCases::ConstantValuedVariables(Int32).0.flag2\ := False;
                        \ConstantsUsingCases::ConstantValuedVariables(Int32).0.num6\ := to_signed(163, 32);
                        \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State\ := \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_4\ => 
                        -- True branch of the if-else started in state \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_2\.
                        \ConstantsUsingCases::ConstantValuedVariables(Int32).0.num5\ := to_signed(13, 32);
                        -- Going to the state after the if-else which was started in state \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_2\.
                        if (\ConstantsUsingCases::ConstantValuedVariables(Int32).0._State\ = \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_4\) then 
                            \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State\ := \ConstantsUsingCases::ConstantValuedVariables(Int32).0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases::ConstantValuedVariables(System.Int32).0 state machine end


    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases::ConstantPassingToMethod(System.Int32).0 state machine start
    \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._StateMachine\: process (\Clock\) 
        Variable \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._State\: \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._States\ := \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._State_0\;
        Variable \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.input\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.num\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.num2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.num3\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.return.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.binaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._Finished\ <= false;
                \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).input1.parameter.Out.0\ <= to_signed(0, 32);
                \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).input2.parameter.Out.0\ <= to_signed(0, 32);
                \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.ConstantsUsingCases::ConstantUsingMethod(Int32,Int32)._Started.0\ <= false;
                \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._State\ := \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._State_0\;
                \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.input\ := to_signed(0, 32);
                \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.num\ := to_signed(0, 32);
                \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.num2\ := to_signed(0, 32);
                \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.num3\ := to_signed(0, 32);
                \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.return.0\ := to_signed(0, 32);
                \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.binaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._State\ is 
                    when \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ConstantsUsingCases::ConstantPassingToMethod(Int32).0._Started\ = true) then 
                            \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._State\ := \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ConstantsUsingCases::ConstantPassingToMethod(Int32).0._Started\ = true) then 
                            \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._Finished\ <= true;
                        else 
                            \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._Finished\ <= false;
                            \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._State\ := \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._State_2\ => 
                        \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.input\ := \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.input.parameter.In\;
                        \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.num\ := to_signed(15, 32);
                        \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.num2\ := to_signed(145, 32);
                        -- Starting state machine invocation for the following method: System.Int32 Hast.TestInputs.Various.ConstantsUsingCases::ConstantUsingMethod(System.Int32,System.Int32)
                        \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).input1.parameter.Out.0\ <= to_signed(145, 32);
                        \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).input2.parameter.Out.0\ <= \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.input\;
                        \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.ConstantsUsingCases::ConstantUsingMethod(Int32,Int32)._Started.0\ <= true;
                        \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._State\ := \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Int32 Hast.TestInputs.Various.ConstantsUsingCases::ConstantUsingMethod(System.Int32,System.Int32)
                        if (\ConstantsUsingCases::ConstantPassingToMethod(Int32).0.ConstantsUsingCases::ConstantUsingMethod(Int32,Int32)._Started.0\ = \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.ConstantsUsingCases::ConstantUsingMethod(Int32,Int32)._Finished.0\) then 
                            \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.ConstantsUsingCases::ConstantUsingMethod(Int32,Int32)._Started.0\ <= false;
                            \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.return.0\ := \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).return.0\;
                            \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.binaryOperationResult.0\ := \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.return.0\ + to_signed(298, 32);
                            \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.num3\ := \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.binaryOperationResult.0\;
                            \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._State\ := \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases::ConstantPassingToMethod(System.Int32).0 state machine end


    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases::ConstantPassingToObject().0 state machine start
    \ConstantsUsingCases::ConstantPassingToObject().0._StateMachine\: process (\Clock\) 
        Variable \ConstantsUsingCases::ConstantPassingToObject().0._State\: \ConstantsUsingCases::ConstantPassingToObject().0._States\ := \ConstantsUsingCases::ConstantPassingToObject().0._State_0\;
        Variable \ConstantsUsingCases::ConstantPassingToObject().0.num\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ConstantsUsingCases::ConstantPassingToObject().0.array\: \unsigned32_Array\(0 to 4) := (others => to_unsigned(0, 32));
        Variable \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
        Variable \ConstantsUsingCases::ConstantPassingToObject().0.array2\: \unsigned32_Array\(0 to 4) := (others => to_unsigned(0, 32));
        Variable \ConstantsUsingCases::ConstantPassingToObject().0.arrayLength\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ConstantsUsingCases::ConstantPassingToObject().0.arrayLengthCopy\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ConstantsUsingCases::ConstantPassingToObject().0.nonSubstitutableArrayLengthCopy\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder2\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
        Variable \ConstantsUsingCases::ConstantPassingToObject().0.previous\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
        Variable \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder3\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
        Variable \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder4\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
        Variable \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder5\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1\;
        Variable \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder6\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder2\;
        Variable \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder7\: \Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder2\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ConstantsUsingCases::ConstantPassingToObject().0._Finished\ <= false;
                \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).array.parameter.Out.0\ <= (others => to_unsigned(0, 32));
                \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Started.0\ <= false;
                \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).size.parameter.Out.0\ <= to_unsigned(0, 32);
                \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32)._Started.0\ <= false;
                \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1)._Started.0\ <= false;
                \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).size.parameter.Out.0\ <= to_unsigned(0, 32);
                \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32)._Started.0\ <= false;
                \ConstantsUsingCases::ConstantPassingToObject().0._State\ := \ConstantsUsingCases::ConstantPassingToObject().0._State_0\;
                \ConstantsUsingCases::ConstantPassingToObject().0.num\ := to_signed(0, 32);
                \ConstantsUsingCases::ConstantPassingToObject().0.array\ := (others => to_unsigned(0, 32));
                \ConstantsUsingCases::ConstantPassingToObject().0.array2\ := (others => to_unsigned(0, 32));
                \ConstantsUsingCases::ConstantPassingToObject().0.arrayLength\ := to_unsigned(0, 32);
                \ConstantsUsingCases::ConstantPassingToObject().0.arrayLengthCopy\ := to_unsigned(0, 32);
                \ConstantsUsingCases::ConstantPassingToObject().0.nonSubstitutableArrayLengthCopy\ := to_unsigned(0, 32);
            else 
                case \ConstantsUsingCases::ConstantPassingToObject().0._State\ is 
                    when \ConstantsUsingCases::ConstantPassingToObject().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ConstantsUsingCases::ConstantPassingToObject().0._Started\ = true) then 
                            \ConstantsUsingCases::ConstantPassingToObject().0._State\ := \ConstantsUsingCases::ConstantPassingToObject().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases::ConstantPassingToObject().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ConstantsUsingCases::ConstantPassingToObject().0._Started\ = true) then 
                            \ConstantsUsingCases::ConstantPassingToObject().0._Finished\ <= true;
                        else 
                            \ConstantsUsingCases::ConstantPassingToObject().0._Finished\ <= false;
                            \ConstantsUsingCases::ConstantPassingToObject().0._State\ := \ConstantsUsingCases::ConstantPassingToObject().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases::ConstantPassingToObject().0._State_2\ => 
                        \ConstantsUsingCases::ConstantPassingToObject().0.num\ := to_signed(5, 32);
                        \ConstantsUsingCases::ConstantPassingToObject().0.array\ := (others => to_unsigned(0, 32));
                        -- Initializing record fields to their defaults.
                        \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder\.\IsNull\ := false;
                        \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder\.\ArrayLength\ := to_unsigned(0, 32);
                        \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder\.\ArrayLengthCopy\ := to_unsigned(0, 32);
                        \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder\.\NonSubstitutableArrayLengthCopy\ := to_unsigned(0, 32);
                        \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder\.\Array\ := (others => to_unsigned(0, 32));
                        -- Invoking the target's constructor.
                        -- Starting state machine invocation for the following method: System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32[])
                        \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).this.parameter.Out.0\ <= \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder\;
                        \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).array.parameter.Out.0\ <= \ConstantsUsingCases::ConstantPassingToObject().0.array\;
                        \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Started.0\ <= true;
                        \ConstantsUsingCases::ConstantPassingToObject().0._State\ := \ConstantsUsingCases::ConstantPassingToObject().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases::ConstantPassingToObject().0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32[])
                        if (\ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Started.0\ = \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Finished.0\) then 
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Started.0\ <= false;
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder\ := \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).this.parameter.In.0\;
                            \ConstantsUsingCases::ConstantPassingToObject().0.array\ := \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).array.parameter.In.0\;
                            \ConstantsUsingCases::ConstantPassingToObject().0.array2\ := \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder\.\Array\;
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayLength\ := to_unsigned(5, 32);
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayLengthCopy\ := to_unsigned(160, 32);
                            \ConstantsUsingCases::ConstantPassingToObject().0.nonSubstitutableArrayLengthCopy\ := \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder\.\NonSubstitutableArrayLengthCopy\;
                            -- Initializing record fields to their defaults.
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder2\.\IsNull\ := false;
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder2\.\ArrayLength\ := to_unsigned(0, 32);
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder2\.\ArrayLengthCopy\ := to_unsigned(0, 32);
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder2\.\NonSubstitutableArrayLengthCopy\ := to_unsigned(0, 32);
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder2\.\Array\ := (others => to_unsigned(0, 32));
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32[])
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).this.parameter.Out.0\ <= \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder2\;
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).array.parameter.Out.0\ <= \ConstantsUsingCases::ConstantPassingToObject().0.array2\;
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Started.0\ <= true;
                            \ConstantsUsingCases::ConstantPassingToObject().0._State\ := \ConstantsUsingCases::ConstantPassingToObject().0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases::ConstantPassingToObject().0._State_4\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32[])
                        if (\ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Started.0\ = \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Finished.0\) then 
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Started.0\ <= false;
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder2\ := \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).this.parameter.In.0\;
                            \ConstantsUsingCases::ConstantPassingToObject().0.array2\ := \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).array.parameter.In.0\;
                            -- Initializing record fields to their defaults.
                            \ConstantsUsingCases::ConstantPassingToObject().0.previous\.\IsNull\ := false;
                            \ConstantsUsingCases::ConstantPassingToObject().0.previous\.\ArrayLength\ := to_unsigned(0, 32);
                            \ConstantsUsingCases::ConstantPassingToObject().0.previous\.\ArrayLengthCopy\ := to_unsigned(0, 32);
                            \ConstantsUsingCases::ConstantPassingToObject().0.previous\.\NonSubstitutableArrayLengthCopy\ := to_unsigned(0, 32);
                            \ConstantsUsingCases::ConstantPassingToObject().0.previous\.\Array\ := (others => to_unsigned(0, 32));
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32)
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).this.parameter.Out.0\ <= \ConstantsUsingCases::ConstantPassingToObject().0.previous\;
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).size.parameter.Out.0\ <= to_unsigned(5, 32);
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32)._Started.0\ <= true;
                            \ConstantsUsingCases::ConstantPassingToObject().0._State\ := \ConstantsUsingCases::ConstantPassingToObject().0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases::ConstantPassingToObject().0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32)
                        if (\ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32)._Started.0\ = \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32)._Finished.0\) then 
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32)._Started.0\ <= false;
                            \ConstantsUsingCases::ConstantPassingToObject().0.previous\ := \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).this.parameter.In.0\;
                            -- Initializing record fields to their defaults.
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder3\.\IsNull\ := false;
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder3\.\ArrayLength\ := to_unsigned(0, 32);
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder3\.\ArrayLengthCopy\ := to_unsigned(0, 32);
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder3\.\NonSubstitutableArrayLengthCopy\ := to_unsigned(0, 32);
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder3\.\Array\ := (others => to_unsigned(0, 32));
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32)
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).this.parameter.Out.0\ <= \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder3\;
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).size.parameter.Out.0\ <= to_unsigned(5, 32);
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32)._Started.0\ <= true;
                            \ConstantsUsingCases::ConstantPassingToObject().0._State\ := \ConstantsUsingCases::ConstantPassingToObject().0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases::ConstantPassingToObject().0._State_6\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32)
                        if (\ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32)._Started.0\ = \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32)._Finished.0\) then 
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32)._Started.0\ <= false;
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder3\ := \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).this.parameter.In.0\;
                            -- Initializing record fields to their defaults.
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder4\.\IsNull\ := false;
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder4\.\ArrayLength\ := to_unsigned(0, 32);
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder4\.\ArrayLengthCopy\ := to_unsigned(0, 32);
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder4\.\NonSubstitutableArrayLengthCopy\ := to_unsigned(0, 32);
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder4\.\Array\ := (others => to_unsigned(0, 32));
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32)
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).this.parameter.Out.0\ <= \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder4\;
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).size.parameter.Out.0\ <= to_unsigned(5, 32);
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32)._Started.0\ <= true;
                            \ConstantsUsingCases::ConstantPassingToObject().0._State\ := \ConstantsUsingCases::ConstantPassingToObject().0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases::ConstantPassingToObject().0._State_7\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32)
                        if (\ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32)._Started.0\ = \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32)._Finished.0\) then 
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32)._Started.0\ <= false;
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder4\ := \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).this.parameter.In.0\;
                            -- Initializing record fields to their defaults.
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder5\.\IsNull\ := false;
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder5\.\ArrayLength\ := to_unsigned(0, 32);
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder5\.\ArrayLengthCopy\ := to_unsigned(0, 32);
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder5\.\NonSubstitutableArrayLengthCopy\ := to_unsigned(0, 32);
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder5\.\Array\ := (others => to_unsigned(0, 32));
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1)
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).this.parameter.Out.0\ <= \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder5\;
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).previous.parameter.Out.0\ <= \ConstantsUsingCases::ConstantPassingToObject().0.previous\;
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1)._Started.0\ <= true;
                            \ConstantsUsingCases::ConstantPassingToObject().0._State\ := \ConstantsUsingCases::ConstantPassingToObject().0._State_8\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases::ConstantPassingToObject().0._State_8\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1)
                        if (\ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1)._Started.0\ = \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1)._Finished.0\) then 
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1)._Started.0\ <= false;
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder5\ := \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).this.parameter.In.0\;
                            \ConstantsUsingCases::ConstantPassingToObject().0.previous\ := \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).previous.parameter.In.0\;
                            -- Initializing record fields to their defaults.
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder6\.\IsNull\ := false;
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder6\.\ArrayLength\ := to_unsigned(0, 32);
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder2::.ctor(System.UInt32)
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).this.parameter.Out.0\ <= \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder6\;
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).size.parameter.Out.0\ <= to_unsigned(5, 32);
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32)._Started.0\ <= true;
                            \ConstantsUsingCases::ConstantPassingToObject().0._State\ := \ConstantsUsingCases::ConstantPassingToObject().0._State_9\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases::ConstantPassingToObject().0._State_9\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder2::.ctor(System.UInt32)
                        if (\ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32)._Started.0\ = \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32)._Finished.0\) then 
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32)._Started.0\ <= false;
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder6\ := \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).this.parameter.In.0\;
                            -- Initializing record fields to their defaults.
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder7\.\IsNull\ := false;
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder7\.\ArrayLength\ := to_unsigned(0, 32);
                            -- Invoking the target's constructor.
                            -- Starting state machine invocation for the following method: System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder2::.ctor(System.UInt32)
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).this.parameter.Out.0\ <= \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder7\;
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).size.parameter.Out.0\ <= to_unsigned(13, 32);
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32)._Started.0\ <= true;
                            \ConstantsUsingCases::ConstantPassingToObject().0._State\ := \ConstantsUsingCases::ConstantPassingToObject().0._State_10\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases::ConstantPassingToObject().0._State_10\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder2::.ctor(System.UInt32)
                        if (\ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32)._Started.0\ = \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32)._Finished.0\) then 
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32)._Started.0\ <= false;
                            \ConstantsUsingCases::ConstantPassingToObject().0.arrayHolder7\ := \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).this.parameter.In.0\;
                            \ConstantsUsingCases::ConstantPassingToObject().0._State\ := \ConstantsUsingCases::ConstantPassingToObject().0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.Various.ConstantsUsingCases::ConstantPassingToObject().0 state machine end


    -- System.Int32 Hast.TestInputs.Various.ConstantsUsingCases::ConstantUsingMethod(System.Int32,System.Int32).0 state machine start
    \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._StateMachine\: process (\Clock\) 
        Variable \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._State\: \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._States\ := \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._State_0\;
        Variable \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0.input1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0.input2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0.binaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._Finished\ <= false;
                \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0.return\ <= to_signed(0, 32);
                \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._State\ := \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._State_0\;
                \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0.input1\ := to_signed(0, 32);
                \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0.input2\ := to_signed(0, 32);
                \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0.binaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._State\ is 
                    when \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._Started\ = true) then 
                            \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._State\ := \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._Started\ = true) then 
                            \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._Finished\ <= true;
                        else 
                            \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._Finished\ <= false;
                            \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._State\ := \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._State_2\ => 
                        \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0.input1\ := \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0.input1.parameter.In\;
                        \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0.input2\ := \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0.input2.parameter.In\;
                        \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0.binaryOperationResult.0\ := to_signed(298, 32) - \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0.input2\;
                        \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0.return\ <= \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0.binaryOperationResult.0\;
                        \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._State\ := \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.Int32 Hast.TestInputs.Various.ConstantsUsingCases::ConstantUsingMethod(System.Int32,System.Int32).0 state machine end


    -- System.Void Hast.TestInputs.Various.LoopCases::BreakInLoop(System.Int32).0 state machine start
    \LoopCases::BreakInLoop(Int32).0._StateMachine\: process (\Clock\) 
        Variable \LoopCases::BreakInLoop(Int32).0._State\: \LoopCases::BreakInLoop(Int32).0._States\ := \LoopCases::BreakInLoop(Int32).0._State_0\;
        Variable \LoopCases::BreakInLoop(Int32).0.input\: signed(31 downto 0) := to_signed(0, 32);
        Variable \LoopCases::BreakInLoop(Int32).0.num\: signed(31 downto 0) := to_signed(0, 32);
        Variable \LoopCases::BreakInLoop(Int32).0.i\: signed(31 downto 0) := to_signed(0, 32);
        Variable \LoopCases::BreakInLoop(Int32).0.flag\: boolean := false;
        Variable \LoopCases::BreakInLoop(Int32).0.binaryOperationResult.0\: boolean := false;
        Variable \LoopCases::BreakInLoop(Int32).0.binaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \LoopCases::BreakInLoop(Int32).0.binaryOperationResult.2\: boolean := false;
        Variable \LoopCases::BreakInLoop(Int32).0.binaryOperationResult.3\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \LoopCases::BreakInLoop(Int32).0._Finished\ <= false;
                \LoopCases::BreakInLoop(Int32).0._State\ := \LoopCases::BreakInLoop(Int32).0._State_0\;
                \LoopCases::BreakInLoop(Int32).0.input\ := to_signed(0, 32);
                \LoopCases::BreakInLoop(Int32).0.num\ := to_signed(0, 32);
                \LoopCases::BreakInLoop(Int32).0.i\ := to_signed(0, 32);
                \LoopCases::BreakInLoop(Int32).0.flag\ := false;
                \LoopCases::BreakInLoop(Int32).0.binaryOperationResult.0\ := false;
                \LoopCases::BreakInLoop(Int32).0.binaryOperationResult.1\ := to_signed(0, 32);
                \LoopCases::BreakInLoop(Int32).0.binaryOperationResult.2\ := false;
                \LoopCases::BreakInLoop(Int32).0.binaryOperationResult.3\ := to_signed(0, 32);
            else 
                case \LoopCases::BreakInLoop(Int32).0._State\ is 
                    when \LoopCases::BreakInLoop(Int32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\LoopCases::BreakInLoop(Int32).0._Started\ = true) then 
                            \LoopCases::BreakInLoop(Int32).0._State\ := \LoopCases::BreakInLoop(Int32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \LoopCases::BreakInLoop(Int32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\LoopCases::BreakInLoop(Int32).0._Started\ = true) then 
                            \LoopCases::BreakInLoop(Int32).0._Finished\ <= true;
                        else 
                            \LoopCases::BreakInLoop(Int32).0._Finished\ <= false;
                            \LoopCases::BreakInLoop(Int32).0._State\ := \LoopCases::BreakInLoop(Int32).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \LoopCases::BreakInLoop(Int32).0._State_2\ => 
                        \LoopCases::BreakInLoop(Int32).0.input\ := \LoopCases::BreakInLoop(Int32).0.input.parameter.In\;
                        \LoopCases::BreakInLoop(Int32).0.num\ := \LoopCases::BreakInLoop(Int32).0.input\;
                        \LoopCases::BreakInLoop(Int32).0.i\ := to_signed(0, 32);
                        -- Starting a while loop.
                        \LoopCases::BreakInLoop(Int32).0._State\ := \LoopCases::BreakInLoop(Int32).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \LoopCases::BreakInLoop(Int32).0._State_3\ => 
                        -- Repeated state of the while loop which was started in state \LoopCases::BreakInLoop(Int32).0._State_2\.
                        -- The while loop's condition:
                        \LoopCases::BreakInLoop(Int32).0.binaryOperationResult.0\ := \LoopCases::BreakInLoop(Int32).0.i\ < \LoopCases::BreakInLoop(Int32).0.input\;
                        if (\LoopCases::BreakInLoop(Int32).0.binaryOperationResult.0\) then 
                            \LoopCases::BreakInLoop(Int32).0.binaryOperationResult.1\ := \LoopCases::BreakInLoop(Int32).0.num\ + \LoopCases::BreakInLoop(Int32).0.i\;
                            \LoopCases::BreakInLoop(Int32).0.num\ := \LoopCases::BreakInLoop(Int32).0.binaryOperationResult.1\;
                            \LoopCases::BreakInLoop(Int32).0.binaryOperationResult.2\ := \LoopCases::BreakInLoop(Int32).0.num\ > to_signed(10, 32);
                            \LoopCases::BreakInLoop(Int32).0.flag\ := \LoopCases::BreakInLoop(Int32).0.binaryOperationResult.2\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \LoopCases::BreakInLoop(Int32).0._State_6\ and ends in state \LoopCases::BreakInLoop(Int32).0._State_6\.
                            --     * Execution after either branch will continue in the following state: \LoopCases::BreakInLoop(Int32).0._State_5\.

                            if (\LoopCases::BreakInLoop(Int32).0.flag\) then 
                                \LoopCases::BreakInLoop(Int32).0._State\ := \LoopCases::BreakInLoop(Int32).0._State_6\;
                            else 
                                -- There was no false branch, so going directly to the state after the if-else.
                                \LoopCases::BreakInLoop(Int32).0._State\ := \LoopCases::BreakInLoop(Int32).0._State_5\;
                            end if;
                        else 
                            \LoopCases::BreakInLoop(Int32).0._State\ := \LoopCases::BreakInLoop(Int32).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \LoopCases::BreakInLoop(Int32).0._State_4\ => 
                        -- State after the while loop which was started in state \LoopCases::BreakInLoop(Int32).0._State_2\.
                        \LoopCases::BreakInLoop(Int32).0._State\ := \LoopCases::BreakInLoop(Int32).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \LoopCases::BreakInLoop(Int32).0._State_5\ => 
                        -- State after the if-else which was started in state \LoopCases::BreakInLoop(Int32).0._State_3\.
                        \LoopCases::BreakInLoop(Int32).0.binaryOperationResult.3\ := \LoopCases::BreakInLoop(Int32).0.i\ + to_signed(1, 32);
                        \LoopCases::BreakInLoop(Int32).0.i\ := \LoopCases::BreakInLoop(Int32).0.binaryOperationResult.3\;
                        -- Returning to the repeated state of the while loop which was started in state \LoopCases::BreakInLoop(Int32).0._State_2\ if the loop wasn't exited with a state change.
                        if (\LoopCases::BreakInLoop(Int32).0._State\ = \LoopCases::BreakInLoop(Int32).0._State_5\) then 
                            \LoopCases::BreakInLoop(Int32).0._State\ := \LoopCases::BreakInLoop(Int32).0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \LoopCases::BreakInLoop(Int32).0._State_6\ => 
                        -- True branch of the if-else started in state \LoopCases::BreakInLoop(Int32).0._State_3\.
                        -- Exiting the while loop with a break statement.
                        \LoopCases::BreakInLoop(Int32).0._State\ := \LoopCases::BreakInLoop(Int32).0._State_4\;
                        -- Going to the state after the if-else which was started in state \LoopCases::BreakInLoop(Int32).0._State_3\.
                        if (\LoopCases::BreakInLoop(Int32).0._State\ = \LoopCases::BreakInLoop(Int32).0._State_6\) then 
                            \LoopCases::BreakInLoop(Int32).0._State\ := \LoopCases::BreakInLoop(Int32).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.Various.LoopCases::BreakInLoop(System.Int32).0 state machine end


    -- System.Void Hast.TestInputs.Various.LoopCases::BreakInLoopInLoop(System.Int32).0 state machine start
    \LoopCases::BreakInLoopInLoop(Int32).0._StateMachine\: process (\Clock\) 
        Variable \LoopCases::BreakInLoopInLoop(Int32).0._State\: \LoopCases::BreakInLoopInLoop(Int32).0._States\ := \LoopCases::BreakInLoopInLoop(Int32).0._State_0\;
        Variable \LoopCases::BreakInLoopInLoop(Int32).0.input\: signed(31 downto 0) := to_signed(0, 32);
        Variable \LoopCases::BreakInLoopInLoop(Int32).0.num\: signed(31 downto 0) := to_signed(0, 32);
        Variable \LoopCases::BreakInLoopInLoop(Int32).0.i\: signed(31 downto 0) := to_signed(0, 32);
        Variable \LoopCases::BreakInLoopInLoop(Int32).0.j\: signed(31 downto 0) := to_signed(0, 32);
        Variable \LoopCases::BreakInLoopInLoop(Int32).0.flag\: boolean := false;
        Variable \LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.0\: boolean := false;
        Variable \LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.1\: boolean := false;
        Variable \LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.3\: boolean := false;
        Variable \LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.4\: signed(31 downto 0) := to_signed(0, 32);
        Variable \LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.5\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \LoopCases::BreakInLoopInLoop(Int32).0._Finished\ <= false;
                \LoopCases::BreakInLoopInLoop(Int32).0._State\ := \LoopCases::BreakInLoopInLoop(Int32).0._State_0\;
                \LoopCases::BreakInLoopInLoop(Int32).0.input\ := to_signed(0, 32);
                \LoopCases::BreakInLoopInLoop(Int32).0.num\ := to_signed(0, 32);
                \LoopCases::BreakInLoopInLoop(Int32).0.i\ := to_signed(0, 32);
                \LoopCases::BreakInLoopInLoop(Int32).0.j\ := to_signed(0, 32);
                \LoopCases::BreakInLoopInLoop(Int32).0.flag\ := false;
                \LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.0\ := false;
                \LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.1\ := false;
                \LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.2\ := to_signed(0, 32);
                \LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.3\ := false;
                \LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.4\ := to_signed(0, 32);
                \LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.5\ := to_signed(0, 32);
            else 
                case \LoopCases::BreakInLoopInLoop(Int32).0._State\ is 
                    when \LoopCases::BreakInLoopInLoop(Int32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\LoopCases::BreakInLoopInLoop(Int32).0._Started\ = true) then 
                            \LoopCases::BreakInLoopInLoop(Int32).0._State\ := \LoopCases::BreakInLoopInLoop(Int32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \LoopCases::BreakInLoopInLoop(Int32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\LoopCases::BreakInLoopInLoop(Int32).0._Started\ = true) then 
                            \LoopCases::BreakInLoopInLoop(Int32).0._Finished\ <= true;
                        else 
                            \LoopCases::BreakInLoopInLoop(Int32).0._Finished\ <= false;
                            \LoopCases::BreakInLoopInLoop(Int32).0._State\ := \LoopCases::BreakInLoopInLoop(Int32).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \LoopCases::BreakInLoopInLoop(Int32).0._State_2\ => 
                        \LoopCases::BreakInLoopInLoop(Int32).0.input\ := \LoopCases::BreakInLoopInLoop(Int32).0.input.parameter.In\;
                        \LoopCases::BreakInLoopInLoop(Int32).0.num\ := \LoopCases::BreakInLoopInLoop(Int32).0.input\;
                        \LoopCases::BreakInLoopInLoop(Int32).0.i\ := to_signed(0, 32);
                        -- Starting a while loop.
                        \LoopCases::BreakInLoopInLoop(Int32).0._State\ := \LoopCases::BreakInLoopInLoop(Int32).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \LoopCases::BreakInLoopInLoop(Int32).0._State_3\ => 
                        -- Repeated state of the while loop which was started in state \LoopCases::BreakInLoopInLoop(Int32).0._State_2\.
                        -- The while loop's condition:
                        \LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.0\ := \LoopCases::BreakInLoopInLoop(Int32).0.i\ < \LoopCases::BreakInLoopInLoop(Int32).0.input\;
                        if (\LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.0\) then 
                            \LoopCases::BreakInLoopInLoop(Int32).0.j\ := to_signed(0, 32);
                            -- Starting a while loop.
                            \LoopCases::BreakInLoopInLoop(Int32).0._State\ := \LoopCases::BreakInLoopInLoop(Int32).0._State_5\;
                        else 
                            \LoopCases::BreakInLoopInLoop(Int32).0._State\ := \LoopCases::BreakInLoopInLoop(Int32).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \LoopCases::BreakInLoopInLoop(Int32).0._State_4\ => 
                        -- State after the while loop which was started in state \LoopCases::BreakInLoopInLoop(Int32).0._State_2\.
                        \LoopCases::BreakInLoopInLoop(Int32).0._State\ := \LoopCases::BreakInLoopInLoop(Int32).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \LoopCases::BreakInLoopInLoop(Int32).0._State_5\ => 
                        -- Repeated state of the while loop which was started in state \LoopCases::BreakInLoopInLoop(Int32).0._State_3\.
                        -- The while loop's condition:
                        \LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.1\ := \LoopCases::BreakInLoopInLoop(Int32).0.j\ < \LoopCases::BreakInLoopInLoop(Int32).0.i\;
                        if (\LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.1\) then 
                            \LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.2\ := \LoopCases::BreakInLoopInLoop(Int32).0.num\ + \LoopCases::BreakInLoopInLoop(Int32).0.i\;
                            \LoopCases::BreakInLoopInLoop(Int32).0.num\ := \LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.2\;
                            \LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.3\ := \LoopCases::BreakInLoopInLoop(Int32).0.num\ > to_signed(10, 32);
                            \LoopCases::BreakInLoopInLoop(Int32).0.flag\ := \LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.3\;

                            -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                            --     * The true branch starts in state \LoopCases::BreakInLoopInLoop(Int32).0._State_8\ and ends in state \LoopCases::BreakInLoopInLoop(Int32).0._State_8\.
                            --     * Execution after either branch will continue in the following state: \LoopCases::BreakInLoopInLoop(Int32).0._State_7\.

                            if (\LoopCases::BreakInLoopInLoop(Int32).0.flag\) then 
                                \LoopCases::BreakInLoopInLoop(Int32).0._State\ := \LoopCases::BreakInLoopInLoop(Int32).0._State_8\;
                            else 
                                -- There was no false branch, so going directly to the state after the if-else.
                                \LoopCases::BreakInLoopInLoop(Int32).0._State\ := \LoopCases::BreakInLoopInLoop(Int32).0._State_7\;
                            end if;
                        else 
                            \LoopCases::BreakInLoopInLoop(Int32).0._State\ := \LoopCases::BreakInLoopInLoop(Int32).0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.3
                    when \LoopCases::BreakInLoopInLoop(Int32).0._State_6\ => 
                        -- State after the while loop which was started in state \LoopCases::BreakInLoopInLoop(Int32).0._State_3\.
                        \LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.5\ := \LoopCases::BreakInLoopInLoop(Int32).0.i\ + to_signed(1, 32);
                        \LoopCases::BreakInLoopInLoop(Int32).0.i\ := \LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.5\;
                        -- Returning to the repeated state of the while loop which was started in state \LoopCases::BreakInLoopInLoop(Int32).0._State_2\ if the loop wasn't exited with a state change.
                        if (\LoopCases::BreakInLoopInLoop(Int32).0._State\ = \LoopCases::BreakInLoopInLoop(Int32).0._State_6\) then 
                            \LoopCases::BreakInLoopInLoop(Int32).0._State\ := \LoopCases::BreakInLoopInLoop(Int32).0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \LoopCases::BreakInLoopInLoop(Int32).0._State_7\ => 
                        -- State after the if-else which was started in state \LoopCases::BreakInLoopInLoop(Int32).0._State_5\.
                        \LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.4\ := \LoopCases::BreakInLoopInLoop(Int32).0.j\ + to_signed(1, 32);
                        \LoopCases::BreakInLoopInLoop(Int32).0.j\ := \LoopCases::BreakInLoopInLoop(Int32).0.binaryOperationResult.4\;
                        -- Returning to the repeated state of the while loop which was started in state \LoopCases::BreakInLoopInLoop(Int32).0._State_3\ if the loop wasn't exited with a state change.
                        if (\LoopCases::BreakInLoopInLoop(Int32).0._State\ = \LoopCases::BreakInLoopInLoop(Int32).0._State_7\) then 
                            \LoopCases::BreakInLoopInLoop(Int32).0._State\ := \LoopCases::BreakInLoopInLoop(Int32).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \LoopCases::BreakInLoopInLoop(Int32).0._State_8\ => 
                        -- True branch of the if-else started in state \LoopCases::BreakInLoopInLoop(Int32).0._State_5\.
                        -- Exiting the while loop with a break statement.
                        \LoopCases::BreakInLoopInLoop(Int32).0._State\ := \LoopCases::BreakInLoopInLoop(Int32).0._State_6\;
                        -- Going to the state after the if-else which was started in state \LoopCases::BreakInLoopInLoop(Int32).0._State_5\.
                        if (\LoopCases::BreakInLoopInLoop(Int32).0._State\ = \LoopCases::BreakInLoopInLoop(Int32).0._State_8\) then 
                            \LoopCases::BreakInLoopInLoop(Int32).0._State\ := \LoopCases::BreakInLoopInLoop(Int32).0._State_7\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.Various.LoopCases::BreakInLoopInLoop(System.Int32).0 state machine end


    -- System.Void Hast.TestInputs.Various.ObjectUsingCases::NullUsage().0 state machine start
    \ObjectUsingCases::NullUsage().0._StateMachine\: process (\Clock\) 
        Variable \ObjectUsingCases::NullUsage().0._State\: \ObjectUsingCases::NullUsage().0._States\ := \ObjectUsingCases::NullUsage().0._State_0\;
        Variable \ObjectUsingCases::NullUsage().0.myClass\: \Hast.TestInputs.Various.ObjectUsingCases/MyClass\;
        Variable \ObjectUsingCases::NullUsage().0.flag\: boolean := false;
        Variable \ObjectUsingCases::NullUsage().0.flag2\: boolean := false;
        Variable \ObjectUsingCases::NullUsage().0.binaryOperationResult.0\: boolean := false;
        Variable \ObjectUsingCases::NullUsage().0.binaryOperationResult.1\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ObjectUsingCases::NullUsage().0._Finished\ <= false;
                \ObjectUsingCases::NullUsage().0._State\ := \ObjectUsingCases::NullUsage().0._State_0\;
                \ObjectUsingCases::NullUsage().0.flag\ := false;
                \ObjectUsingCases::NullUsage().0.flag2\ := false;
                \ObjectUsingCases::NullUsage().0.binaryOperationResult.0\ := false;
                \ObjectUsingCases::NullUsage().0.binaryOperationResult.1\ := false;
            else 
                case \ObjectUsingCases::NullUsage().0._State\ is 
                    when \ObjectUsingCases::NullUsage().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ObjectUsingCases::NullUsage().0._Started\ = true) then 
                            \ObjectUsingCases::NullUsage().0._State\ := \ObjectUsingCases::NullUsage().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectUsingCases::NullUsage().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ObjectUsingCases::NullUsage().0._Started\ = true) then 
                            \ObjectUsingCases::NullUsage().0._Finished\ <= true;
                        else 
                            \ObjectUsingCases::NullUsage().0._Finished\ <= false;
                            \ObjectUsingCases::NullUsage().0._State\ := \ObjectUsingCases::NullUsage().0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectUsingCases::NullUsage().0._State_2\ => 
                        -- Initializing record fields to their defaults.
                        \ObjectUsingCases::NullUsage().0.myClass\.\IsNull\ := false;
                        \ObjectUsingCases::NullUsage().0.myClass\.\MyProperty\ := to_signed(0, 32);
                        \ObjectUsingCases::NullUsage().0.myClass\.\MyProperty\ := to_signed(5, 32);
                        \ObjectUsingCases::NullUsage().0.binaryOperationResult.0\ := \ObjectUsingCases::NullUsage().0.myClass\.\IsNull\ = true;
                        \ObjectUsingCases::NullUsage().0.flag\ := \ObjectUsingCases::NullUsage().0.binaryOperationResult.0\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \ObjectUsingCases::NullUsage().0._State_4\ and ends in state \ObjectUsingCases::NullUsage().0._State_4\.
                        --     * Execution after either branch will continue in the following state: \ObjectUsingCases::NullUsage().0._State_3\.

                        if (\ObjectUsingCases::NullUsage().0.flag\) then 
                            \ObjectUsingCases::NullUsage().0._State\ := \ObjectUsingCases::NullUsage().0._State_4\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \ObjectUsingCases::NullUsage().0._State\ := \ObjectUsingCases::NullUsage().0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ObjectUsingCases::NullUsage().0._State_3\ => 
                        -- State after the if-else which was started in state \ObjectUsingCases::NullUsage().0._State_2\.
                        \ObjectUsingCases::NullUsage().0.myClass\.\IsNull\ := true;
                        \ObjectUsingCases::NullUsage().0.binaryOperationResult.1\ := \ObjectUsingCases::NullUsage().0.myClass\.\IsNull\ /= true;
                        \ObjectUsingCases::NullUsage().0.flag2\ := \ObjectUsingCases::NullUsage().0.binaryOperationResult.1\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \ObjectUsingCases::NullUsage().0._State_6\ and ends in state \ObjectUsingCases::NullUsage().0._State_6\.
                        --     * Execution after either branch will continue in the following state: \ObjectUsingCases::NullUsage().0._State_5\.

                        if (\ObjectUsingCases::NullUsage().0.flag2\) then 
                            \ObjectUsingCases::NullUsage().0._State\ := \ObjectUsingCases::NullUsage().0._State_6\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \ObjectUsingCases::NullUsage().0._State\ := \ObjectUsingCases::NullUsage().0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ObjectUsingCases::NullUsage().0._State_4\ => 
                        -- True branch of the if-else started in state \ObjectUsingCases::NullUsage().0._State_2\.
                        -- Initializing record fields to their defaults.
                        \ObjectUsingCases::NullUsage().0.myClass\.\IsNull\ := false;
                        \ObjectUsingCases::NullUsage().0.myClass\.\MyProperty\ := to_signed(0, 32);
                        -- Going to the state after the if-else which was started in state \ObjectUsingCases::NullUsage().0._State_2\.
                        if (\ObjectUsingCases::NullUsage().0._State\ = \ObjectUsingCases::NullUsage().0._State_4\) then 
                            \ObjectUsingCases::NullUsage().0._State\ := \ObjectUsingCases::NullUsage().0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectUsingCases::NullUsage().0._State_5\ => 
                        -- State after the if-else which was started in state \ObjectUsingCases::NullUsage().0._State_3\.
                        \ObjectUsingCases::NullUsage().0._State\ := \ObjectUsingCases::NullUsage().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectUsingCases::NullUsage().0._State_6\ => 
                        -- True branch of the if-else started in state \ObjectUsingCases::NullUsage().0._State_3\.
                        \ObjectUsingCases::NullUsage().0.myClass\.\MyProperty\ := to_signed(10, 32);
                        -- Going to the state after the if-else which was started in state \ObjectUsingCases::NullUsage().0._State_3\.
                        if (\ObjectUsingCases::NullUsage().0._State\ = \ObjectUsingCases::NullUsage().0._State_6\) then 
                            \ObjectUsingCases::NullUsage().0._State\ := \ObjectUsingCases::NullUsage().0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.Various.ObjectUsingCases::NullUsage().0 state machine end


    -- System.Void Hast.TestInputs.Various.ObjectUsingCases::VoidReturn(System.Int32).0 state machine start
    \ObjectUsingCases::VoidReturn(Int32).0._StateMachine\: process (\Clock\) 
        Variable \ObjectUsingCases::VoidReturn(Int32).0._State\: \ObjectUsingCases::VoidReturn(Int32).0._States\ := \ObjectUsingCases::VoidReturn(Int32).0._State_0\;
        Variable \ObjectUsingCases::VoidReturn(Int32).0.input\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ObjectUsingCases::VoidReturn(Int32).0.myClass\: \Hast.TestInputs.Various.ObjectUsingCases/MyClass\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ObjectUsingCases::VoidReturn(Int32).0._Finished\ <= false;
                \ObjectUsingCases::VoidReturn(Int32).0.ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass)._Started.0\ <= false;
                \ObjectUsingCases::VoidReturn(Int32).0._State\ := \ObjectUsingCases::VoidReturn(Int32).0._State_0\;
                \ObjectUsingCases::VoidReturn(Int32).0.input\ := to_signed(0, 32);
            else 
                case \ObjectUsingCases::VoidReturn(Int32).0._State\ is 
                    when \ObjectUsingCases::VoidReturn(Int32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ObjectUsingCases::VoidReturn(Int32).0._Started\ = true) then 
                            \ObjectUsingCases::VoidReturn(Int32).0._State\ := \ObjectUsingCases::VoidReturn(Int32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectUsingCases::VoidReturn(Int32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ObjectUsingCases::VoidReturn(Int32).0._Started\ = true) then 
                            \ObjectUsingCases::VoidReturn(Int32).0._Finished\ <= true;
                        else 
                            \ObjectUsingCases::VoidReturn(Int32).0._Finished\ <= false;
                            \ObjectUsingCases::VoidReturn(Int32).0._State\ := \ObjectUsingCases::VoidReturn(Int32).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectUsingCases::VoidReturn(Int32).0._State_2\ => 
                        \ObjectUsingCases::VoidReturn(Int32).0.input\ := \ObjectUsingCases::VoidReturn(Int32).0.input.parameter.In\;
                        -- Initializing record fields to their defaults.
                        \ObjectUsingCases::VoidReturn(Int32).0.myClass\.\IsNull\ := false;
                        \ObjectUsingCases::VoidReturn(Int32).0.myClass\.\MyProperty\ := to_signed(0, 32);
                        \ObjectUsingCases::VoidReturn(Int32).0.myClass\.\MyProperty\ := \ObjectUsingCases::VoidReturn(Int32).0.input\;
                        -- Starting state machine invocation for the following method: System.Void Hast.TestInputs.Various.ObjectUsingCases::VoidMethod(Hast.TestInputs.Various.ObjectUsingCases/MyClass)
                        \ObjectUsingCases::VoidReturn(Int32).0.ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).myClass.parameter.Out.0\ <= \ObjectUsingCases::VoidReturn(Int32).0.myClass\;
                        \ObjectUsingCases::VoidReturn(Int32).0.ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass)._Started.0\ <= true;
                        \ObjectUsingCases::VoidReturn(Int32).0._State\ := \ObjectUsingCases::VoidReturn(Int32).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectUsingCases::VoidReturn(Int32).0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Void Hast.TestInputs.Various.ObjectUsingCases::VoidMethod(Hast.TestInputs.Various.ObjectUsingCases/MyClass)
                        if (\ObjectUsingCases::VoidReturn(Int32).0.ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass)._Started.0\ = \ObjectUsingCases::VoidReturn(Int32).0.ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass)._Finished.0\) then 
                            \ObjectUsingCases::VoidReturn(Int32).0.ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass)._Started.0\ <= false;
                            \ObjectUsingCases::VoidReturn(Int32).0.myClass\ := \ObjectUsingCases::VoidReturn(Int32).0.ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).myClass.parameter.In.0\;
                            \ObjectUsingCases::VoidReturn(Int32).0._State\ := \ObjectUsingCases::VoidReturn(Int32).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.Various.ObjectUsingCases::VoidReturn(System.Int32).0 state machine end


    -- System.Void Hast.TestInputs.Various.ObjectUsingCases::VoidMethod(Hast.TestInputs.Various.ObjectUsingCases/MyClass).0 state machine start
    \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._StateMachine\: process (\Clock\) 
        Variable \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State\: \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._States\ := \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_0\;
        Variable \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.myClass\: \Hast.TestInputs.Various.ObjectUsingCases/MyClass\;
        Variable \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.flag\: boolean := false;
        Variable \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.flag2\: boolean := false;
        Variable \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.binaryOperationResult.0\: boolean := false;
        Variable \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.binaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.binaryOperationResult.2\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._Finished\ <= false;
                \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State\ := \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_0\;
                \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.flag\ := false;
                \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.flag2\ := false;
                \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.binaryOperationResult.0\ := false;
                \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.binaryOperationResult.1\ := to_signed(0, 32);
                \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.binaryOperationResult.2\ := false;
            else 
                case \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State\ is 
                    when \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._Started\ = true) then 
                            \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State\ := \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._Started\ = true) then 
                            \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._Finished\ <= true;
                        else 
                            \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._Finished\ <= false;
                            \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State\ := \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.myClass.parameter.Out\ <= \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.myClass\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_2\ => 
                        \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.myClass\ := \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.myClass.parameter.In\;
                        \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.binaryOperationResult.0\ := \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.myClass\.\MyProperty\ < to_signed(10, 32);
                        \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.flag\ := \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.binaryOperationResult.0\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_4\ and ends in state \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_5\.
                        --     * Execution after either branch will continue in the following state: \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_3\.

                        if (\ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.flag\) then 
                            \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State\ := \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_4\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State\ := \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_3\ => 
                        -- State after the if-else which was started in state \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_2\.
                        \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.myClass\.\MyProperty\ := to_signed(5, 32);
                        \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State\ := \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_4\ => 
                        -- True branch of the if-else started in state \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_2\.
                        \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.binaryOperationResult.1\ := resize(\ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.myClass\.\MyProperty\ * to_signed(10, 32), 32);
                        \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.myClass\.\MyProperty\ := \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.binaryOperationResult.1\;
                        \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.binaryOperationResult.2\ := \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.myClass\.\MyProperty\ = to_signed(10, 32);
                        \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.flag2\ := \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.binaryOperationResult.2\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_6\ and ends in state \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_6\.
                        --     * Execution after either branch will continue in the following state: \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_5\.

                        if (\ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.flag2\) then 
                            \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State\ := \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_6\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State\ := \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_5\ => 
                        -- State after the if-else which was started in state \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_4\.
                        -- Going to the state after the if-else which was started in state \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_2\.
                        if (\ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State\ = \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_5\) then 
                            \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State\ := \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_6\ => 
                        -- True branch of the if-else started in state \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_4\.
                        \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State\ := \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_1\;
                        -- Going to the state after the if-else which was started in state \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_4\.
                        if (\ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State\ = \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_6\) then 
                            \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State\ := \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._State_5\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.Various.ObjectUsingCases::VoidMethod(Hast.TestInputs.Various.ObjectUsingCases/MyClass).0 state machine end


    -- System.Boolean Hast.TestInputs.Various.ParallelCases/Calculator::IsEven().0 state machine start
    \ParallelCases/Calculator::IsEven().0._StateMachine\: process (\Clock\) 
        Variable \ParallelCases/Calculator::IsEven().0._State\: \ParallelCases/Calculator::IsEven().0._States\ := \ParallelCases/Calculator::IsEven().0._State_0\;
        Variable \ParallelCases/Calculator::IsEven().0.this\: \Hast.TestInputs.Various.ParallelCases/Calculator\;
        Variable \ParallelCases/Calculator::IsEven().0.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/Calculator::IsEven().0.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ParallelCases/Calculator::IsEven().0.binaryOperationResult.1\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ParallelCases/Calculator::IsEven().0._Finished\ <= false;
                \ParallelCases/Calculator::IsEven().0.return\ <= false;
                \ParallelCases/Calculator::IsEven().0._State\ := \ParallelCases/Calculator::IsEven().0._State_0\;
                \ParallelCases/Calculator::IsEven().0.binaryOperationResult.0\ := to_unsigned(0, 32);
                \ParallelCases/Calculator::IsEven().0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                \ParallelCases/Calculator::IsEven().0.binaryOperationResult.1\ := false;
            else 
                case \ParallelCases/Calculator::IsEven().0._State\ is 
                    when \ParallelCases/Calculator::IsEven().0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ParallelCases/Calculator::IsEven().0._Started\ = true) then 
                            \ParallelCases/Calculator::IsEven().0._State\ := \ParallelCases/Calculator::IsEven().0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases/Calculator::IsEven().0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ParallelCases/Calculator::IsEven().0._Started\ = true) then 
                            \ParallelCases/Calculator::IsEven().0._Finished\ <= true;
                        else 
                            \ParallelCases/Calculator::IsEven().0._Finished\ <= false;
                            \ParallelCases/Calculator::IsEven().0._State\ := \ParallelCases/Calculator::IsEven().0._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \ParallelCases/Calculator::IsEven().0.this.parameter.Out\ <= \ParallelCases/Calculator::IsEven().0.this\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases/Calculator::IsEven().0._State_2\ => 
                        \ParallelCases/Calculator::IsEven().0.this\ := \ParallelCases/Calculator::IsEven().0.this.parameter.In\;
                        \ParallelCases/Calculator::IsEven().0._State\ := \ParallelCases/Calculator::IsEven().0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases/Calculator::IsEven().0._State_3\ => 
                        -- Waiting for the result to appear in \ParallelCases/Calculator::IsEven().0.binaryOperationResult.0\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\ParallelCases/Calculator::IsEven().0.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \ParallelCases/Calculator::IsEven().0._State\ := \ParallelCases/Calculator::IsEven().0._State_4\;
                            \ParallelCases/Calculator::IsEven().0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \ParallelCases/Calculator::IsEven().0.clockCyclesWaitedForBinaryOperationResult.0\ := \ParallelCases/Calculator::IsEven().0.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        \ParallelCases/Calculator::IsEven().0.binaryOperationResult.0\ := \ParallelCases/Calculator::IsEven().0.this\.\Number\ mod to_unsigned(2, 32);
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \ParallelCases/Calculator::IsEven().0._State_4\ => 
                        \ParallelCases/Calculator::IsEven().0.binaryOperationResult.1\ := \ParallelCases/Calculator::IsEven().0.binaryOperationResult.0\ = to_unsigned(0, 32);
                        \ParallelCases/Calculator::IsEven().0.return\ <= \ParallelCases/Calculator::IsEven().0.binaryOperationResult.1\;
                        \ParallelCases/Calculator::IsEven().0._State\ := \ParallelCases/Calculator::IsEven().0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.TestInputs.Various.ParallelCases/Calculator::IsEven().0 state machine end


    -- System.Boolean Hast.TestInputs.Various.ParallelCases/Calculator::IsEven().1 state machine start
    \ParallelCases/Calculator::IsEven().1._StateMachine\: process (\Clock\) 
        Variable \ParallelCases/Calculator::IsEven().1._State\: \ParallelCases/Calculator::IsEven().1._States\ := \ParallelCases/Calculator::IsEven().1._State_0\;
        Variable \ParallelCases/Calculator::IsEven().1.this\: \Hast.TestInputs.Various.ParallelCases/Calculator\;
        Variable \ParallelCases/Calculator::IsEven().1.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/Calculator::IsEven().1.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ParallelCases/Calculator::IsEven().1.binaryOperationResult.1\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ParallelCases/Calculator::IsEven().1._Finished\ <= false;
                \ParallelCases/Calculator::IsEven().1.return\ <= false;
                \ParallelCases/Calculator::IsEven().1._State\ := \ParallelCases/Calculator::IsEven().1._State_0\;
                \ParallelCases/Calculator::IsEven().1.binaryOperationResult.0\ := to_unsigned(0, 32);
                \ParallelCases/Calculator::IsEven().1.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                \ParallelCases/Calculator::IsEven().1.binaryOperationResult.1\ := false;
            else 
                case \ParallelCases/Calculator::IsEven().1._State\ is 
                    when \ParallelCases/Calculator::IsEven().1._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ParallelCases/Calculator::IsEven().1._Started\ = true) then 
                            \ParallelCases/Calculator::IsEven().1._State\ := \ParallelCases/Calculator::IsEven().1._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases/Calculator::IsEven().1._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ParallelCases/Calculator::IsEven().1._Started\ = true) then 
                            \ParallelCases/Calculator::IsEven().1._Finished\ <= true;
                        else 
                            \ParallelCases/Calculator::IsEven().1._Finished\ <= false;
                            \ParallelCases/Calculator::IsEven().1._State\ := \ParallelCases/Calculator::IsEven().1._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \ParallelCases/Calculator::IsEven().1.this.parameter.Out\ <= \ParallelCases/Calculator::IsEven().1.this\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases/Calculator::IsEven().1._State_2\ => 
                        \ParallelCases/Calculator::IsEven().1.this\ := \ParallelCases/Calculator::IsEven().1.this.parameter.In\;
                        \ParallelCases/Calculator::IsEven().1._State\ := \ParallelCases/Calculator::IsEven().1._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases/Calculator::IsEven().1._State_3\ => 
                        -- Waiting for the result to appear in \ParallelCases/Calculator::IsEven().1.binaryOperationResult.0\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\ParallelCases/Calculator::IsEven().1.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \ParallelCases/Calculator::IsEven().1._State\ := \ParallelCases/Calculator::IsEven().1._State_4\;
                            \ParallelCases/Calculator::IsEven().1.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \ParallelCases/Calculator::IsEven().1.clockCyclesWaitedForBinaryOperationResult.0\ := \ParallelCases/Calculator::IsEven().1.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        \ParallelCases/Calculator::IsEven().1.binaryOperationResult.0\ := \ParallelCases/Calculator::IsEven().1.this\.\Number\ mod to_unsigned(2, 32);
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \ParallelCases/Calculator::IsEven().1._State_4\ => 
                        \ParallelCases/Calculator::IsEven().1.binaryOperationResult.1\ := \ParallelCases/Calculator::IsEven().1.binaryOperationResult.0\ = to_unsigned(0, 32);
                        \ParallelCases/Calculator::IsEven().1.return\ <= \ParallelCases/Calculator::IsEven().1.binaryOperationResult.1\;
                        \ParallelCases/Calculator::IsEven().1._State\ := \ParallelCases/Calculator::IsEven().1._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.TestInputs.Various.ParallelCases/Calculator::IsEven().1 state machine end


    -- System.Boolean Hast.TestInputs.Various.ParallelCases/Calculator::IsEven().2 state machine start
    \ParallelCases/Calculator::IsEven().2._StateMachine\: process (\Clock\) 
        Variable \ParallelCases/Calculator::IsEven().2._State\: \ParallelCases/Calculator::IsEven().2._States\ := \ParallelCases/Calculator::IsEven().2._State_0\;
        Variable \ParallelCases/Calculator::IsEven().2.this\: \Hast.TestInputs.Various.ParallelCases/Calculator\;
        Variable \ParallelCases/Calculator::IsEven().2.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/Calculator::IsEven().2.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ParallelCases/Calculator::IsEven().2.binaryOperationResult.1\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ParallelCases/Calculator::IsEven().2._Finished\ <= false;
                \ParallelCases/Calculator::IsEven().2.return\ <= false;
                \ParallelCases/Calculator::IsEven().2._State\ := \ParallelCases/Calculator::IsEven().2._State_0\;
                \ParallelCases/Calculator::IsEven().2.binaryOperationResult.0\ := to_unsigned(0, 32);
                \ParallelCases/Calculator::IsEven().2.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                \ParallelCases/Calculator::IsEven().2.binaryOperationResult.1\ := false;
            else 
                case \ParallelCases/Calculator::IsEven().2._State\ is 
                    when \ParallelCases/Calculator::IsEven().2._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ParallelCases/Calculator::IsEven().2._Started\ = true) then 
                            \ParallelCases/Calculator::IsEven().2._State\ := \ParallelCases/Calculator::IsEven().2._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases/Calculator::IsEven().2._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ParallelCases/Calculator::IsEven().2._Started\ = true) then 
                            \ParallelCases/Calculator::IsEven().2._Finished\ <= true;
                        else 
                            \ParallelCases/Calculator::IsEven().2._Finished\ <= false;
                            \ParallelCases/Calculator::IsEven().2._State\ := \ParallelCases/Calculator::IsEven().2._State_0\;
                        end if;
                        -- Writing back out-flowing parameters so any changes made in this state machine will be reflected in the invoking one too.
                        \ParallelCases/Calculator::IsEven().2.this.parameter.Out\ <= \ParallelCases/Calculator::IsEven().2.this\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases/Calculator::IsEven().2._State_2\ => 
                        \ParallelCases/Calculator::IsEven().2.this\ := \ParallelCases/Calculator::IsEven().2.this.parameter.In\;
                        \ParallelCases/Calculator::IsEven().2._State\ := \ParallelCases/Calculator::IsEven().2._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases/Calculator::IsEven().2._State_3\ => 
                        -- Waiting for the result to appear in \ParallelCases/Calculator::IsEven().2.binaryOperationResult.0\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\ParallelCases/Calculator::IsEven().2.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \ParallelCases/Calculator::IsEven().2._State\ := \ParallelCases/Calculator::IsEven().2._State_4\;
                            \ParallelCases/Calculator::IsEven().2.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \ParallelCases/Calculator::IsEven().2.clockCyclesWaitedForBinaryOperationResult.0\ := \ParallelCases/Calculator::IsEven().2.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        \ParallelCases/Calculator::IsEven().2.binaryOperationResult.0\ := \ParallelCases/Calculator::IsEven().2.this\.\Number\ mod to_unsigned(2, 32);
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \ParallelCases/Calculator::IsEven().2._State_4\ => 
                        \ParallelCases/Calculator::IsEven().2.binaryOperationResult.1\ := \ParallelCases/Calculator::IsEven().2.binaryOperationResult.0\ = to_unsigned(0, 32);
                        \ParallelCases/Calculator::IsEven().2.return\ <= \ParallelCases/Calculator::IsEven().2.binaryOperationResult.1\;
                        \ParallelCases/Calculator::IsEven().2._State\ := \ParallelCases/Calculator::IsEven().2._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.TestInputs.Various.ParallelCases/Calculator::IsEven().2 state machine end


    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(System.UInt32).0 state machine start
    \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._StateMachine\: process (\Clock\) 
        Variable \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State\: \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._States\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State_0\;
        Variable \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.indexObject\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.binaryOperationResult.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.binaryOperationResult.2\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._Finished\ <= false;
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.return\ <= false;
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State_0\;
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.indexObject\ := to_unsigned(0, 32);
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.num\ := to_unsigned(0, 32);
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.binaryOperationResult.0\ := to_unsigned(0, 32);
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.binaryOperationResult.1\ := to_unsigned(0, 32);
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.binaryOperationResult.2\ := false;
            else 
                case \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State\ is 
                    when \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._Started\ = true) then 
                            \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._Started\ = true) then 
                            \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._Finished\ <= true;
                        else 
                            \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._Finished\ <= false;
                            \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State_2\ => 
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.indexObject\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.indexObject.parameter.In\;
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.num\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.indexObject\;
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.binaryOperationResult.0\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.num\ + \System.UInt32 Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::input\;
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.num\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.binaryOperationResult.0\;
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State_3\ => 
                        -- Waiting for the result to appear in \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.binaryOperationResult.1\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State_4\;
                            \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.binaryOperationResult.1\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.num\ mod to_unsigned(2, 32);
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State_4\ => 
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.binaryOperationResult.2\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.binaryOperationResult.1\ = to_unsigned(0, 32);
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.return\ <= \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.binaryOperationResult.2\;
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(System.UInt32).0 state machine end


    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(System.UInt32).1 state machine start
    \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._StateMachine\: process (\Clock\) 
        Variable \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State\: \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._States\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State_0\;
        Variable \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.indexObject\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.binaryOperationResult.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.binaryOperationResult.2\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._Finished\ <= false;
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.return\ <= false;
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State_0\;
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.indexObject\ := to_unsigned(0, 32);
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.num\ := to_unsigned(0, 32);
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.binaryOperationResult.0\ := to_unsigned(0, 32);
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.binaryOperationResult.1\ := to_unsigned(0, 32);
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.binaryOperationResult.2\ := false;
            else 
                case \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State\ is 
                    when \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._Started\ = true) then 
                            \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._Started\ = true) then 
                            \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._Finished\ <= true;
                        else 
                            \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._Finished\ <= false;
                            \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State_2\ => 
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.indexObject\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.indexObject.parameter.In\;
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.num\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.indexObject\;
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.binaryOperationResult.0\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.num\ + \System.UInt32 Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::input\;
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.num\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.binaryOperationResult.0\;
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State_3\ => 
                        -- Waiting for the result to appear in \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.binaryOperationResult.1\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State_4\;
                            \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.clockCyclesWaitedForBinaryOperationResult.0\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.binaryOperationResult.1\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.num\ mod to_unsigned(2, 32);
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State_4\ => 
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.binaryOperationResult.2\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.binaryOperationResult.1\ = to_unsigned(0, 32);
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.return\ <= \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.binaryOperationResult.2\;
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(System.UInt32).1 state machine end


    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(System.UInt32).2 state machine start
    \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._StateMachine\: process (\Clock\) 
        Variable \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State\: \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._States\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State_0\;
        Variable \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.indexObject\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.binaryOperationResult.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.binaryOperationResult.2\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._Finished\ <= false;
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.return\ <= false;
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State_0\;
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.indexObject\ := to_unsigned(0, 32);
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.num\ := to_unsigned(0, 32);
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.binaryOperationResult.0\ := to_unsigned(0, 32);
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.binaryOperationResult.1\ := to_unsigned(0, 32);
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.binaryOperationResult.2\ := false;
            else 
                case \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State\ is 
                    when \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._Started\ = true) then 
                            \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._Started\ = true) then 
                            \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._Finished\ <= true;
                        else 
                            \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._Finished\ <= false;
                            \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State_2\ => 
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.indexObject\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.indexObject.parameter.In\;
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.num\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.indexObject\;
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.binaryOperationResult.0\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.num\ + \System.UInt32 Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::input\;
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.num\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.binaryOperationResult.0\;
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State_3\ => 
                        -- Waiting for the result to appear in \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.binaryOperationResult.1\ (have to wait 7 clock cycles in this state).
                        -- The assignment needs to be kept up for multi-cycle operations for the result to actually appear in the target.
                        if (\ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(7, 32)) then 
                            \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State_4\;
                            \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.clockCyclesWaitedForBinaryOperationResult.0\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.binaryOperationResult.1\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.num\ mod to_unsigned(2, 32);
                        -- Clock cycles needed to complete this state (approximation): 7
                    when \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State_4\ => 
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.binaryOperationResult.2\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.binaryOperationResult.1\ = to_unsigned(0, 32);
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.return\ <= \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.binaryOperationResult.2\;
                        \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State\ := \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(System.UInt32).2 state machine end


    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(System.UInt32).0 state machine start
    \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._StateMachine\: process (\Clock\) 
        Variable \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._State\: \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._States\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._State_0\;
        Variable \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.indexObject\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.objectdc3e2eea384e7e52700cea72b1c1cb21eb3ce1928d378edcac638af24735332f\: \Hast.TestInputs.Various.ParallelCases/Calculator\;
        Variable \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.return.0\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._Finished\ <= false;
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.return\ <= false;
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.ParallelCases/Calculator::IsEven()._Started.0\ <= false;
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._State\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._State_0\;
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.indexObject\ := to_unsigned(0, 32);
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.num\ := to_unsigned(0, 32);
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.binaryOperationResult.0\ := to_unsigned(0, 32);
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.return.0\ := false;
            else 
                case \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._State\ is 
                    when \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._Started\ = true) then 
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._State\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._Started\ = true) then 
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._Finished\ <= true;
                        else 
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._Finished\ <= false;
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._State\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._State_2\ => 
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.indexObject\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.indexObject.parameter.In\;
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.num\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.indexObject\;
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.binaryOperationResult.0\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.num\ + \System.UInt32 Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::input\;
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.num\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.binaryOperationResult.0\;
                        -- Initializing record fields to their defaults.
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.objectdc3e2eea384e7e52700cea72b1c1cb21eb3ce1928d378edcac638af24735332f\.\IsNull\ := false;
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.objectdc3e2eea384e7e52700cea72b1c1cb21eb3ce1928d378edcac638af24735332f\.\Number\ := to_unsigned(0, 32);
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.objectdc3e2eea384e7e52700cea72b1c1cb21eb3ce1928d378edcac638af24735332f\.\Number\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.num\;
                        -- Starting state machine invocation for the following method: System.Boolean Hast.TestInputs.Various.ParallelCases/Calculator::IsEven()
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.ParallelCases/Calculator::IsEven().this.parameter.Out.0\ <= \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.objectdc3e2eea384e7e52700cea72b1c1cb21eb3ce1928d378edcac638af24735332f\;
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.ParallelCases/Calculator::IsEven()._Started.0\ <= true;
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._State\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Hast.TestInputs.Various.ParallelCases/Calculator::IsEven()
                        if (\ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.ParallelCases/Calculator::IsEven()._Started.0\ = \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.ParallelCases/Calculator::IsEven()._Finished.0\) then 
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.ParallelCases/Calculator::IsEven()._Started.0\ <= false;
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.return.0\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.ParallelCases/Calculator::IsEven().return.0\;
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.objectdc3e2eea384e7e52700cea72b1c1cb21eb3ce1928d378edcac638af24735332f\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.ParallelCases/Calculator::IsEven().this.parameter.In.0\;
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.return\ <= \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.return.0\;
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._State\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(System.UInt32).0 state machine end


    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(System.UInt32).1 state machine start
    \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._StateMachine\: process (\Clock\) 
        Variable \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._State\: \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._States\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._State_0\;
        Variable \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.indexObject\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.objectdc3e2eea384e7e52700cea72b1c1cb21eb3ce1928d378edcac638af24735332f\: \Hast.TestInputs.Various.ParallelCases/Calculator\;
        Variable \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.return.0\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._Finished\ <= false;
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.return\ <= false;
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.ParallelCases/Calculator::IsEven()._Started.0\ <= false;
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._State\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._State_0\;
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.indexObject\ := to_unsigned(0, 32);
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.num\ := to_unsigned(0, 32);
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.binaryOperationResult.0\ := to_unsigned(0, 32);
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.return.0\ := false;
            else 
                case \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._State\ is 
                    when \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._Started\ = true) then 
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._State\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._Started\ = true) then 
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._Finished\ <= true;
                        else 
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._Finished\ <= false;
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._State\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._State_2\ => 
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.indexObject\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.indexObject.parameter.In\;
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.num\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.indexObject\;
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.binaryOperationResult.0\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.num\ + \System.UInt32 Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::input\;
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.num\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.binaryOperationResult.0\;
                        -- Initializing record fields to their defaults.
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.objectdc3e2eea384e7e52700cea72b1c1cb21eb3ce1928d378edcac638af24735332f\.\IsNull\ := false;
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.objectdc3e2eea384e7e52700cea72b1c1cb21eb3ce1928d378edcac638af24735332f\.\Number\ := to_unsigned(0, 32);
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.objectdc3e2eea384e7e52700cea72b1c1cb21eb3ce1928d378edcac638af24735332f\.\Number\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.num\;
                        -- Starting state machine invocation for the following method: System.Boolean Hast.TestInputs.Various.ParallelCases/Calculator::IsEven()
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.ParallelCases/Calculator::IsEven().this.parameter.Out.0\ <= \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.objectdc3e2eea384e7e52700cea72b1c1cb21eb3ce1928d378edcac638af24735332f\;
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.ParallelCases/Calculator::IsEven()._Started.0\ <= true;
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._State\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Hast.TestInputs.Various.ParallelCases/Calculator::IsEven()
                        if (\ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.ParallelCases/Calculator::IsEven()._Started.0\ = \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.ParallelCases/Calculator::IsEven()._Finished.0\) then 
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.ParallelCases/Calculator::IsEven()._Started.0\ <= false;
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.return.0\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.ParallelCases/Calculator::IsEven().return.0\;
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.objectdc3e2eea384e7e52700cea72b1c1cb21eb3ce1928d378edcac638af24735332f\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.ParallelCases/Calculator::IsEven().this.parameter.In.0\;
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.return\ <= \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.return.0\;
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._State\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(System.UInt32).1 state machine end


    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(System.UInt32).2 state machine start
    \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._StateMachine\: process (\Clock\) 
        Variable \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._State\: \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._States\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._State_0\;
        Variable \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.indexObject\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.objectdc3e2eea384e7e52700cea72b1c1cb21eb3ce1928d378edcac638af24735332f\: \Hast.TestInputs.Various.ParallelCases/Calculator\;
        Variable \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.return.0\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._Finished\ <= false;
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.return\ <= false;
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.ParallelCases/Calculator::IsEven()._Started.0\ <= false;
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._State\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._State_0\;
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.indexObject\ := to_unsigned(0, 32);
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.num\ := to_unsigned(0, 32);
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.binaryOperationResult.0\ := to_unsigned(0, 32);
                \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.return.0\ := false;
            else 
                case \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._State\ is 
                    when \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._Started\ = true) then 
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._State\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._Started\ = true) then 
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._Finished\ <= true;
                        else 
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._Finished\ <= false;
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._State\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._State_2\ => 
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.indexObject\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.indexObject.parameter.In\;
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.num\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.indexObject\;
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.binaryOperationResult.0\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.num\ + \System.UInt32 Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::input\;
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.num\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.binaryOperationResult.0\;
                        -- Initializing record fields to their defaults.
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.objectdc3e2eea384e7e52700cea72b1c1cb21eb3ce1928d378edcac638af24735332f\.\IsNull\ := false;
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.objectdc3e2eea384e7e52700cea72b1c1cb21eb3ce1928d378edcac638af24735332f\.\Number\ := to_unsigned(0, 32);
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.objectdc3e2eea384e7e52700cea72b1c1cb21eb3ce1928d378edcac638af24735332f\.\Number\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.num\;
                        -- Starting state machine invocation for the following method: System.Boolean Hast.TestInputs.Various.ParallelCases/Calculator::IsEven()
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.ParallelCases/Calculator::IsEven().this.parameter.Out.0\ <= \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.objectdc3e2eea384e7e52700cea72b1c1cb21eb3ce1928d378edcac638af24735332f\;
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.ParallelCases/Calculator::IsEven()._Started.0\ <= true;
                        \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._State\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._State_3\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Hast.TestInputs.Various.ParallelCases/Calculator::IsEven()
                        if (\ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.ParallelCases/Calculator::IsEven()._Started.0\ = \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.ParallelCases/Calculator::IsEven()._Finished.0\) then 
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.ParallelCases/Calculator::IsEven()._Started.0\ <= false;
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.return.0\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.ParallelCases/Calculator::IsEven().return.0\;
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.objectdc3e2eea384e7e52700cea72b1c1cb21eb3ce1928d378edcac638af24735332f\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.ParallelCases/Calculator::IsEven().this.parameter.In.0\;
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.return\ <= \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.return.0\;
                            \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._State\ := \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(System.UInt32).2 state machine end


    -- System.Void Hast.TestInputs.Various.ParallelCases::WhenAllWhenAnyAwaitedTasks(System.UInt32).0 state machine start
    \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._StateMachine\: process (\Clock\) 
        Variable \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State\: \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._States\ := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_0\;
        Variable \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.input\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.array\: \boolean_Array\(0 to 2) := (others => false);
        Variable \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.arg_4B_1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.binaryOperationResult.0\: boolean := false;
        Variable \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).invocationIndex\: integer range 0 to 2 := 0;
        Variable \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.binaryOperationResult.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.0\: boolean := false;
        Variable \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.1\: boolean := false;
        Variable \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.2\: boolean := false;
        Variable \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.3\: boolean := false;
        Variable \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.4\: boolean := false;
        Variable \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.5\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._Finished\ <= false;
                \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).indexObject.parameter.Out.0\ <= to_unsigned(0, 32);
                \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.0\ <= false;
                \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).indexObject.parameter.Out.1\ <= to_unsigned(0, 32);
                \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.1\ <= false;
                \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).indexObject.parameter.Out.2\ <= to_unsigned(0, 32);
                \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.2\ <= false;
                \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State\ := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_0\;
                \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.input\ := to_unsigned(0, 32);
                \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.array\ := (others => false);
                \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.num\ := to_unsigned(0, 32);
                \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.arg_4B_1\ := to_signed(0, 32);
                \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.binaryOperationResult.0\ := false;
                \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).invocationIndex\ := 0;
                \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.binaryOperationResult.1\ := to_unsigned(0, 32);
                \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.0\ := false;
                \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.1\ := false;
                \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.2\ := false;
                \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.3\ := false;
                \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.4\ := false;
                \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.5\ := false;
            else 
                case \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State\ is 
                    when \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._Started\ = true) then 
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State\ := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._Started\ = true) then 
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._Finished\ <= true;
                        else 
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._Finished\ <= false;
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State\ := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_2\ => 
                        \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.input\ := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.input.parameter.In\;
                        \System.UInt32 Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::input\ := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.input\;
                        \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.array\ := (others => false);
                        \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.num\ := to_unsigned(0, 32);
                        -- Starting a while loop.
                        \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State\ := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_3\ => 
                        -- Repeated state of the while loop which was started in state \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_2\.
                        -- The while loop's condition:
                        \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.binaryOperationResult.0\ := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.num\ < to_unsigned(3, 32);
                        if (\ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.binaryOperationResult.0\) then 
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.arg_4B_1\ := signed(\ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.num\);
                            -- Starting state machine invocation for the following method: System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(System.UInt32)
                            case \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).invocationIndex\ is 
                                when 0 => 
                                    \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).indexObject.parameter.Out.0\ <= \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.num\;
                                    \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.0\ <= true;
                                when 1 => 
                                    \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).indexObject.parameter.Out.1\ <= \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.num\;
                                    \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.1\ <= true;
                                when 2 => 
                                    \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).indexObject.parameter.Out.2\ <= \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.num\;
                                    \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.2\ <= true;
                            end case;
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).invocationIndex\ := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).invocationIndex\ + 1;
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.binaryOperationResult.1\ := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.num\ + to_unsigned(1, 32);
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.num\ := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.binaryOperationResult.1\;
                        else 
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State\ := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_4\ => 
                        -- State after the while loop which was started in state \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_2\.
                        \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State\ := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_5\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(System.UInt32)
                        if (\ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.1\ = \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Finished.1\ and \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.2\ = \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Finished.2\ and \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.0\ = \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Finished.0\) then 
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.0\ <= false;
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.1\ <= false;
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.2\ <= false;
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).invocationIndex\ := 0;
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.0\ := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).return.0\;
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.1\ := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).return.1\;
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.2\ := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).return.2\;
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.array\(0) := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.0\;
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.array\(1) := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.1\;
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.array\(2) := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.2\;
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State\ := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_6\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_6\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(System.UInt32)
                        if (\ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.1\ = \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Finished.1\ or \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.2\ = \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Finished.2\ or \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.0\ = \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Finished.0\) then 
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.0\ <= false;
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.1\ <= false;
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.2\ <= false;
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).invocationIndex\ := 0;
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.3\ := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).return.0\;
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.4\ := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).return.1\;
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.5\ := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).return.2\;
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.array\(0) := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.3\;
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.array\(1) := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.4\;
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.array\(2) := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.return.5\;
                            \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State\ := \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.Various.ParallelCases::WhenAllWhenAnyAwaitedTasks(System.UInt32).0 state machine end


    -- System.Void Hast.TestInputs.Various.ParallelCases::ObjectUsingTasks(System.UInt32).0 state machine start
    \ParallelCases::ObjectUsingTasks(UInt32).0._StateMachine\: process (\Clock\) 
        Variable \ParallelCases::ObjectUsingTasks(UInt32).0._State\: \ParallelCases::ObjectUsingTasks(UInt32).0._States\ := \ParallelCases::ObjectUsingTasks(UInt32).0._State_0\;
        Variable \ParallelCases::ObjectUsingTasks(UInt32).0.input\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases::ObjectUsingTasks(UInt32).0.array\: \boolean_Array\(0 to 2) := (others => false);
        Variable \ParallelCases::ObjectUsingTasks(UInt32).0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases::ObjectUsingTasks(UInt32).0.arg_4B_1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \ParallelCases::ObjectUsingTasks(UInt32).0.binaryOperationResult.0\: boolean := false;
        Variable \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).invocationIndex\: integer range 0 to 2 := 0;
        Variable \ParallelCases::ObjectUsingTasks(UInt32).0.binaryOperationResult.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \ParallelCases::ObjectUsingTasks(UInt32).0.return.0\: boolean := false;
        Variable \ParallelCases::ObjectUsingTasks(UInt32).0.return.1\: boolean := false;
        Variable \ParallelCases::ObjectUsingTasks(UInt32).0.return.2\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \ParallelCases::ObjectUsingTasks(UInt32).0._Finished\ <= false;
                \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).indexObject.parameter.Out.0\ <= to_unsigned(0, 32);
                \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Started.0\ <= false;
                \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).indexObject.parameter.Out.1\ <= to_unsigned(0, 32);
                \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Started.1\ <= false;
                \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).indexObject.parameter.Out.2\ <= to_unsigned(0, 32);
                \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Started.2\ <= false;
                \ParallelCases::ObjectUsingTasks(UInt32).0._State\ := \ParallelCases::ObjectUsingTasks(UInt32).0._State_0\;
                \ParallelCases::ObjectUsingTasks(UInt32).0.input\ := to_unsigned(0, 32);
                \ParallelCases::ObjectUsingTasks(UInt32).0.array\ := (others => false);
                \ParallelCases::ObjectUsingTasks(UInt32).0.num\ := to_unsigned(0, 32);
                \ParallelCases::ObjectUsingTasks(UInt32).0.arg_4B_1\ := to_signed(0, 32);
                \ParallelCases::ObjectUsingTasks(UInt32).0.binaryOperationResult.0\ := false;
                \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).invocationIndex\ := 0;
                \ParallelCases::ObjectUsingTasks(UInt32).0.binaryOperationResult.1\ := to_unsigned(0, 32);
                \ParallelCases::ObjectUsingTasks(UInt32).0.return.0\ := false;
                \ParallelCases::ObjectUsingTasks(UInt32).0.return.1\ := false;
                \ParallelCases::ObjectUsingTasks(UInt32).0.return.2\ := false;
            else 
                case \ParallelCases::ObjectUsingTasks(UInt32).0._State\ is 
                    when \ParallelCases::ObjectUsingTasks(UInt32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\ParallelCases::ObjectUsingTasks(UInt32).0._Started\ = true) then 
                            \ParallelCases::ObjectUsingTasks(UInt32).0._State\ := \ParallelCases::ObjectUsingTasks(UInt32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases::ObjectUsingTasks(UInt32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\ParallelCases::ObjectUsingTasks(UInt32).0._Started\ = true) then 
                            \ParallelCases::ObjectUsingTasks(UInt32).0._Finished\ <= true;
                        else 
                            \ParallelCases::ObjectUsingTasks(UInt32).0._Finished\ <= false;
                            \ParallelCases::ObjectUsingTasks(UInt32).0._State\ := \ParallelCases::ObjectUsingTasks(UInt32).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases::ObjectUsingTasks(UInt32).0._State_2\ => 
                        \ParallelCases::ObjectUsingTasks(UInt32).0.input\ := \ParallelCases::ObjectUsingTasks(UInt32).0.input.parameter.In\;
                        \System.UInt32 Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::input\ := \ParallelCases::ObjectUsingTasks(UInt32).0.input\;
                        \ParallelCases::ObjectUsingTasks(UInt32).0.array\ := (others => false);
                        \ParallelCases::ObjectUsingTasks(UInt32).0.num\ := to_unsigned(0, 32);
                        -- Starting a while loop.
                        \ParallelCases::ObjectUsingTasks(UInt32).0._State\ := \ParallelCases::ObjectUsingTasks(UInt32).0._State_3\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases::ObjectUsingTasks(UInt32).0._State_3\ => 
                        -- Repeated state of the while loop which was started in state \ParallelCases::ObjectUsingTasks(UInt32).0._State_2\.
                        -- The while loop's condition:
                        \ParallelCases::ObjectUsingTasks(UInt32).0.binaryOperationResult.0\ := \ParallelCases::ObjectUsingTasks(UInt32).0.num\ < to_unsigned(3, 32);
                        if (\ParallelCases::ObjectUsingTasks(UInt32).0.binaryOperationResult.0\) then 
                            \ParallelCases::ObjectUsingTasks(UInt32).0.arg_4B_1\ := signed(\ParallelCases::ObjectUsingTasks(UInt32).0.num\);
                            -- Starting state machine invocation for the following method: System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(System.UInt32)
                            case \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).invocationIndex\ is 
                                when 0 => 
                                    \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).indexObject.parameter.Out.0\ <= \ParallelCases::ObjectUsingTasks(UInt32).0.num\;
                                    \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Started.0\ <= true;
                                when 1 => 
                                    \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).indexObject.parameter.Out.1\ <= \ParallelCases::ObjectUsingTasks(UInt32).0.num\;
                                    \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Started.1\ <= true;
                                when 2 => 
                                    \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).indexObject.parameter.Out.2\ <= \ParallelCases::ObjectUsingTasks(UInt32).0.num\;
                                    \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Started.2\ <= true;
                            end case;
                            \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).invocationIndex\ := \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).invocationIndex\ + 1;
                            \ParallelCases::ObjectUsingTasks(UInt32).0.binaryOperationResult.1\ := \ParallelCases::ObjectUsingTasks(UInt32).0.num\ + to_unsigned(1, 32);
                            \ParallelCases::ObjectUsingTasks(UInt32).0.num\ := \ParallelCases::ObjectUsingTasks(UInt32).0.binaryOperationResult.1\;
                        else 
                            \ParallelCases::ObjectUsingTasks(UInt32).0._State\ := \ParallelCases::ObjectUsingTasks(UInt32).0._State_4\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                    when \ParallelCases::ObjectUsingTasks(UInt32).0._State_4\ => 
                        -- State after the while loop which was started in state \ParallelCases::ObjectUsingTasks(UInt32).0._State_2\.
                        \ParallelCases::ObjectUsingTasks(UInt32).0._State\ := \ParallelCases::ObjectUsingTasks(UInt32).0._State_5\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \ParallelCases::ObjectUsingTasks(UInt32).0._State_5\ => 
                        -- Waiting for the state machine invocation of the following method to finish: System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(System.UInt32)
                        if (\ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Started.1\ = \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Finished.1\ and \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Started.2\ = \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Finished.2\ and \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Started.0\ = \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Finished.0\) then 
                            \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Started.0\ <= false;
                            \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Started.1\ <= false;
                            \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Started.2\ <= false;
                            \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).invocationIndex\ := 0;
                            \ParallelCases::ObjectUsingTasks(UInt32).0.return.0\ := \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).return.0\;
                            \ParallelCases::ObjectUsingTasks(UInt32).0.return.1\ := \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).return.1\;
                            \ParallelCases::ObjectUsingTasks(UInt32).0.return.2\ := \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).return.2\;
                            \ParallelCases::ObjectUsingTasks(UInt32).0.array\(0) := \ParallelCases::ObjectUsingTasks(UInt32).0.return.0\;
                            \ParallelCases::ObjectUsingTasks(UInt32).0.array\(1) := \ParallelCases::ObjectUsingTasks(UInt32).0.return.1\;
                            \ParallelCases::ObjectUsingTasks(UInt32).0.array\(2) := \ParallelCases::ObjectUsingTasks(UInt32).0.return.2\;
                            \ParallelCases::ObjectUsingTasks(UInt32).0._State\ := \ParallelCases::ObjectUsingTasks(UInt32).0._State_1\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.Various.ParallelCases::ObjectUsingTasks(System.UInt32).0 state machine end


    -- System.Void Hast.TestInputs.Various.UnaryCases::IncrementDecrement(System.Int32).0 state machine start
    \UnaryCases::IncrementDecrement(Int32).0._StateMachine\: process (\Clock\) 
        Variable \UnaryCases::IncrementDecrement(Int32).0._State\: \UnaryCases::IncrementDecrement(Int32).0._States\ := \UnaryCases::IncrementDecrement(Int32).0._State_0\;
        Variable \UnaryCases::IncrementDecrement(Int32).0.input\: signed(31 downto 0) := to_signed(0, 32);
        Variable \UnaryCases::IncrementDecrement(Int32).0.array\: \signed32_Array\(0 to 4) := (others => to_signed(0, 32));
        Variable \UnaryCases::IncrementDecrement(Int32).0.flag\: boolean := false;
        Variable \UnaryCases::IncrementDecrement(Int32).0.binaryOperationResult.0\: boolean := false;
        Variable \UnaryCases::IncrementDecrement(Int32).0.binaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \UnaryCases::IncrementDecrement(Int32).0.binaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \UnaryCases::IncrementDecrement(Int32).0._Finished\ <= false;
                \UnaryCases::IncrementDecrement(Int32).0._State\ := \UnaryCases::IncrementDecrement(Int32).0._State_0\;
                \UnaryCases::IncrementDecrement(Int32).0.input\ := to_signed(0, 32);
                \UnaryCases::IncrementDecrement(Int32).0.array\ := (others => to_signed(0, 32));
                \UnaryCases::IncrementDecrement(Int32).0.flag\ := false;
                \UnaryCases::IncrementDecrement(Int32).0.binaryOperationResult.0\ := false;
                \UnaryCases::IncrementDecrement(Int32).0.binaryOperationResult.1\ := to_signed(0, 32);
                \UnaryCases::IncrementDecrement(Int32).0.binaryOperationResult.2\ := to_signed(0, 32);
            else 
                case \UnaryCases::IncrementDecrement(Int32).0._State\ is 
                    when \UnaryCases::IncrementDecrement(Int32).0._State_0\ => 
                        -- Start state
                        -- Waiting for the start signal.
                        if (\UnaryCases::IncrementDecrement(Int32).0._Started\ = true) then 
                            \UnaryCases::IncrementDecrement(Int32).0._State\ := \UnaryCases::IncrementDecrement(Int32).0._State_2\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnaryCases::IncrementDecrement(Int32).0._State_1\ => 
                        -- Final state
                        -- Signaling finished until Started is pulled back to false, then returning to the start state.
                        if (\UnaryCases::IncrementDecrement(Int32).0._Started\ = true) then 
                            \UnaryCases::IncrementDecrement(Int32).0._Finished\ <= true;
                        else 
                            \UnaryCases::IncrementDecrement(Int32).0._Finished\ <= false;
                            \UnaryCases::IncrementDecrement(Int32).0._State\ := \UnaryCases::IncrementDecrement(Int32).0._State_0\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnaryCases::IncrementDecrement(Int32).0._State_2\ => 
                        \UnaryCases::IncrementDecrement(Int32).0.input\ := \UnaryCases::IncrementDecrement(Int32).0.input.parameter.In\;
                        \UnaryCases::IncrementDecrement(Int32).0.array\ := (others => to_signed(0, 32));
                        \UnaryCases::IncrementDecrement(Int32).0.binaryOperationResult.0\ := \UnaryCases::IncrementDecrement(Int32).0.input\ < to_signed(10, 32);
                        \UnaryCases::IncrementDecrement(Int32).0.flag\ := \UnaryCases::IncrementDecrement(Int32).0.binaryOperationResult.0\;

                        -- This if-else was transformed from a .NET if-else. It spans across multiple states:
                        --     * The true branch starts in state \UnaryCases::IncrementDecrement(Int32).0._State_4\ and ends in state \UnaryCases::IncrementDecrement(Int32).0._State_4\.
                        --     * Execution after either branch will continue in the following state: \UnaryCases::IncrementDecrement(Int32).0._State_3\.

                        if (\UnaryCases::IncrementDecrement(Int32).0.flag\) then 
                            \UnaryCases::IncrementDecrement(Int32).0._State\ := \UnaryCases::IncrementDecrement(Int32).0._State_4\;
                        else 
                            -- There was no false branch, so going directly to the state after the if-else.
                            \UnaryCases::IncrementDecrement(Int32).0._State\ := \UnaryCases::IncrementDecrement(Int32).0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.1
                    when \UnaryCases::IncrementDecrement(Int32).0._State_3\ => 
                        -- State after the if-else which was started in state \UnaryCases::IncrementDecrement(Int32).0._State_2\.
                        \UnaryCases::IncrementDecrement(Int32).0._State\ := \UnaryCases::IncrementDecrement(Int32).0._State_1\;
                        -- Clock cycles needed to complete this state (approximation): 0
                    when \UnaryCases::IncrementDecrement(Int32).0._State_4\ => 
                        -- True branch of the if-else started in state \UnaryCases::IncrementDecrement(Int32).0._State_2\.
                        \UnaryCases::IncrementDecrement(Int32).0.array\(to_integer(\UnaryCases::IncrementDecrement(Int32).0.input\)) := to_signed(3, 32);
                        \UnaryCases::IncrementDecrement(Int32).0.binaryOperationResult.1\ := \UnaryCases::IncrementDecrement(Int32).0.input\ + to_signed(1, 32);
                        \UnaryCases::IncrementDecrement(Int32).0.input\ := \UnaryCases::IncrementDecrement(Int32).0.binaryOperationResult.1\;
                        \UnaryCases::IncrementDecrement(Int32).0.array\(to_integer(\UnaryCases::IncrementDecrement(Int32).0.input\)) := to_signed(3, 32);
                        \UnaryCases::IncrementDecrement(Int32).0.binaryOperationResult.2\ := \UnaryCases::IncrementDecrement(Int32).0.input\ - to_signed(1, 32);
                        \UnaryCases::IncrementDecrement(Int32).0.input\ := \UnaryCases::IncrementDecrement(Int32).0.binaryOperationResult.2\;
                        -- Going to the state after the if-else which was started in state \UnaryCases::IncrementDecrement(Int32).0._State_2\.
                        if (\UnaryCases::IncrementDecrement(Int32).0._State\ = \UnaryCases::IncrementDecrement(Int32).0._State_4\) then 
                            \UnaryCases::IncrementDecrement(Int32).0._State\ := \UnaryCases::IncrementDecrement(Int32).0._State_3\;
                        end if;
                        -- Clock cycles needed to complete this state (approximation): 0.2
                end case;
            end if;
        end if;
    end process;
    -- System.Void Hast.TestInputs.Various.UnaryCases::IncrementDecrement(System.Int32).0 state machine end


    -- System.Void Hast::ExternalInvocationProxy() start
    \Finished\ <= \FinishedInternal\;
    \Hast::ExternalInvocationProxy()\: process (\Clock\) 
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \FinishedInternal\ <= false;
                \Hast::ExternalInvocationProxy().RootClass::VirtualMethod(Int32)._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1()._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Interface1Method2()._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Interface2Method1()._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1()._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2()._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::NonVirtualNonInterfaceMehod()._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().StaticClass::StaticMethod()._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().UnusedDeclarations::UnusedMethod()._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().StaticReference::StaticClassUsingMethod()._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().ArrayUsingCases::PassArrayToConstructor()._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().ArrayUsingCases::PassArrayFromMethod()._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().CastingCases::NumberCasting(Int16,Int16)._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantValuedVariables(Int32)._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantPassingToMethod(Int32)._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantPassingToObject()._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().LoopCases::BreakInLoop(Int32)._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().LoopCases::BreakInLoopInLoop(Int32)._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().ObjectUsingCases::NullUsage()._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().ObjectUsingCases::VoidReturn(Int32)._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32)._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().ParallelCases::ObjectUsingTasks(UInt32)._Started.0\ <= false;
                \Hast::ExternalInvocationProxy().UnaryCases::IncrementDecrement(Int32)._Started.0\ <= false;
            else 
                if (\Started\ = true and \FinishedInternal\ = false) then 
                    -- Starting the state machine corresponding to the given member ID.
                    case \MemberId\ is 
                        when 0 => 
                            if (\Hast::ExternalInvocationProxy().RootClass::VirtualMethod(Int32)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().RootClass::VirtualMethod(Int32)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().RootClass::VirtualMethod(Int32)._Started.0\ = \Hast::ExternalInvocationProxy().RootClass::VirtualMethod(Int32)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().RootClass::VirtualMethod(Int32)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 1 => 
                            if (\Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1()._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1()._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1()._Started.0\ = \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1()._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1()._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 2 => 
                            if (\Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Interface1Method2()._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Interface1Method2()._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Interface1Method2()._Started.0\ = \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Interface1Method2()._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Interface1Method2()._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 3 => 
                            if (\Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Interface2Method1()._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Interface2Method1()._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Interface2Method1()._Started.0\ = \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Interface2Method1()._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Interface2Method1()._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 4 => 
                            if (\Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1()._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1()._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1()._Started.0\ = \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1()._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1()._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 5 => 
                            if (\Hast::ExternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2()._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2()._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2()._Started.0\ = \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2()._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2()._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 6 => 
                            if (\Hast::ExternalInvocationProxy().ComplexTypeHierarchy::NonVirtualNonInterfaceMehod()._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::NonVirtualNonInterfaceMehod()._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().ComplexTypeHierarchy::NonVirtualNonInterfaceMehod()._Started.0\ = \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::NonVirtualNonInterfaceMehod()._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::NonVirtualNonInterfaceMehod()._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 7 => 
                            if (\Hast::ExternalInvocationProxy().StaticClass::StaticMethod()._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().StaticClass::StaticMethod()._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().StaticClass::StaticMethod()._Started.0\ = \Hast::ExternalInvocationProxy().StaticClass::StaticMethod()._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().StaticClass::StaticMethod()._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 8 => 
                            if (\Hast::ExternalInvocationProxy().UnusedDeclarations::UnusedMethod()._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().UnusedDeclarations::UnusedMethod()._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().UnusedDeclarations::UnusedMethod()._Started.0\ = \Hast::ExternalInvocationProxy().UnusedDeclarations::UnusedMethod()._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().UnusedDeclarations::UnusedMethod()._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 9 => 
                            if (\Hast::ExternalInvocationProxy().StaticReference::StaticClassUsingMethod()._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().StaticReference::StaticClassUsingMethod()._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().StaticReference::StaticClassUsingMethod()._Started.0\ = \Hast::ExternalInvocationProxy().StaticReference::StaticClassUsingMethod()._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().StaticReference::StaticClassUsingMethod()._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 10 => 
                            if (\Hast::ExternalInvocationProxy().ArrayUsingCases::PassArrayToConstructor()._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().ArrayUsingCases::PassArrayToConstructor()._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().ArrayUsingCases::PassArrayToConstructor()._Started.0\ = \Hast::ExternalInvocationProxy().ArrayUsingCases::PassArrayToConstructor()._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().ArrayUsingCases::PassArrayToConstructor()._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 11 => 
                            if (\Hast::ExternalInvocationProxy().ArrayUsingCases::PassArrayFromMethod()._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().ArrayUsingCases::PassArrayFromMethod()._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().ArrayUsingCases::PassArrayFromMethod()._Started.0\ = \Hast::ExternalInvocationProxy().ArrayUsingCases::PassArrayFromMethod()._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().ArrayUsingCases::PassArrayFromMethod()._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 12 => 
                            if (\Hast::ExternalInvocationProxy().CastingCases::NumberCasting(Int16,Int16)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().CastingCases::NumberCasting(Int16,Int16)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().CastingCases::NumberCasting(Int16,Int16)._Started.0\ = \Hast::ExternalInvocationProxy().CastingCases::NumberCasting(Int16,Int16)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().CastingCases::NumberCasting(Int16,Int16)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 13 => 
                            if (\Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantValuedVariables(Int32)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantValuedVariables(Int32)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantValuedVariables(Int32)._Started.0\ = \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantValuedVariables(Int32)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantValuedVariables(Int32)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 14 => 
                            if (\Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantPassingToMethod(Int32)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantPassingToMethod(Int32)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantPassingToMethod(Int32)._Started.0\ = \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantPassingToMethod(Int32)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantPassingToMethod(Int32)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 15 => 
                            if (\Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantPassingToObject()._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantPassingToObject()._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantPassingToObject()._Started.0\ = \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantPassingToObject()._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantPassingToObject()._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 16 => 
                            if (\Hast::ExternalInvocationProxy().LoopCases::BreakInLoop(Int32)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().LoopCases::BreakInLoop(Int32)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().LoopCases::BreakInLoop(Int32)._Started.0\ = \Hast::ExternalInvocationProxy().LoopCases::BreakInLoop(Int32)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().LoopCases::BreakInLoop(Int32)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 17 => 
                            if (\Hast::ExternalInvocationProxy().LoopCases::BreakInLoopInLoop(Int32)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().LoopCases::BreakInLoopInLoop(Int32)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().LoopCases::BreakInLoopInLoop(Int32)._Started.0\ = \Hast::ExternalInvocationProxy().LoopCases::BreakInLoopInLoop(Int32)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().LoopCases::BreakInLoopInLoop(Int32)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 18 => 
                            if (\Hast::ExternalInvocationProxy().ObjectUsingCases::NullUsage()._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().ObjectUsingCases::NullUsage()._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().ObjectUsingCases::NullUsage()._Started.0\ = \Hast::ExternalInvocationProxy().ObjectUsingCases::NullUsage()._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().ObjectUsingCases::NullUsage()._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 19 => 
                            if (\Hast::ExternalInvocationProxy().ObjectUsingCases::VoidReturn(Int32)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().ObjectUsingCases::VoidReturn(Int32)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().ObjectUsingCases::VoidReturn(Int32)._Started.0\ = \Hast::ExternalInvocationProxy().ObjectUsingCases::VoidReturn(Int32)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().ObjectUsingCases::VoidReturn(Int32)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 20 => 
                            if (\Hast::ExternalInvocationProxy().ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32)._Started.0\ = \Hast::ExternalInvocationProxy().ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 21 => 
                            if (\Hast::ExternalInvocationProxy().ParallelCases::ObjectUsingTasks(UInt32)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().ParallelCases::ObjectUsingTasks(UInt32)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().ParallelCases::ObjectUsingTasks(UInt32)._Started.0\ = \Hast::ExternalInvocationProxy().ParallelCases::ObjectUsingTasks(UInt32)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().ParallelCases::ObjectUsingTasks(UInt32)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when 22 => 
                            if (\Hast::ExternalInvocationProxy().UnaryCases::IncrementDecrement(Int32)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().UnaryCases::IncrementDecrement(Int32)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().UnaryCases::IncrementDecrement(Int32)._Started.0\ = \Hast::ExternalInvocationProxy().UnaryCases::IncrementDecrement(Int32)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().UnaryCases::IncrementDecrement(Int32)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when others => 
                            null;
                    end case;
                else 
                    -- Waiting for Started to be pulled back to zero that signals the framework noting the finish.
                    if (\Started\ = false and \FinishedInternal\ = true) then 
                        \FinishedInternal\ <= false;
                    end if;
                end if;
            end if;
        end if;
    end process;
    -- System.Void Hast::ExternalInvocationProxy() end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::PrivateMethod() start
    \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod()\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::Interface1Method2().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::Interface1Method2().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::Interface1Method2().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::Interface1Method2().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0.runningState.0\ := WaitingForStarted;
                \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0.ComplexTypeHierarchy::PrivateMethod()._Finished.0\ <= false;
                \ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::PrivateMethod()._Finished.0\ <= false;
                \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0.ComplexTypeHierarchy::PrivateMethod()._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0
                case \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0.ComplexTypeHierarchy::PrivateMethod()._Started.0\) then 
                            \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0.ComplexTypeHierarchy::PrivateMethod()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0.runningIndex.0\ := 0;
                            \ComplexTypeHierarchy::PrivateMethod().0._Started\ <= true;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0.runningIndex.0\ is 
                            when 0 => 
                                if (\ComplexTypeHierarchy::PrivateMethod().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0.runningState.0\ := AfterFinished;
                                    \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0.ComplexTypeHierarchy::PrivateMethod()._Finished.0\ <= true;
                                    \ComplexTypeHierarchy::PrivateMethod().0._Started\ <= false;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0.ComplexTypeHierarchy::PrivateMethod()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0.runningState.0\ := WaitingForStarted;
                            \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0.ComplexTypeHierarchy::PrivateMethod()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Interface1Method2().0
                case \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::Interface1Method2().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::PrivateMethod()._Started.0\) then 
                            \ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::PrivateMethod()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::Interface1Method2().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::Interface1Method2().0.runningIndex.0\ := 0;
                            \ComplexTypeHierarchy::PrivateMethod().0._Started\ <= true;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::Interface1Method2().0.runningIndex.0\ is 
                            when 0 => 
                                if (\ComplexTypeHierarchy::PrivateMethod().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::Interface1Method2().0.runningState.0\ := AfterFinished;
                                    \ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::PrivateMethod()._Finished.0\ <= true;
                                    \ComplexTypeHierarchy::PrivateMethod().0._Started\ <= false;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::PrivateMethod()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::Interface1Method2().0.runningState.0\ := WaitingForStarted;
                            \ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::PrivateMethod()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0
                case \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0.ComplexTypeHierarchy::PrivateMethod()._Started.0\) then 
                            \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0.ComplexTypeHierarchy::PrivateMethod()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0.runningIndex.0\ := 0;
                            \ComplexTypeHierarchy::PrivateMethod().0._Started\ <= true;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0.runningIndex.0\ is 
                            when 0 => 
                                if (\ComplexTypeHierarchy::PrivateMethod().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0.runningState.0\ := AfterFinished;
                                    \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0.ComplexTypeHierarchy::PrivateMethod()._Finished.0\ <= true;
                                    \ComplexTypeHierarchy::PrivateMethod().0._Started\ <= false;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0.ComplexTypeHierarchy::PrivateMethod()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::PrivateMethod().ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0.runningState.0\ := WaitingForStarted;
                            \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0.ComplexTypeHierarchy::PrivateMethod()._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::PrivateMethod() end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::StaticMethod() start
    \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod()\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::Interface1Method2().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::Interface1Method2().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::BaseInterfaceMethod2().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::BaseInterfaceMethod2().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::PrivateMethod().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::PrivateMethod().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::Interface1Method2().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::Interface1Method2().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::BaseInterfaceMethod2().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::BaseInterfaceMethod2().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::PrivateMethod().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::PrivateMethod().0.runningState.0\ := WaitingForStarted;
                \ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::StaticMethod()._Finished.0\ <= false;
                \ComplexTypeHierarchy::BaseInterfaceMethod2().0.ComplexTypeHierarchy::StaticMethod()._Finished.0\ <= false;
                \ComplexTypeHierarchy::PrivateMethod().0.ComplexTypeHierarchy::StaticMethod()._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Interface1Method2().0
                case \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::Interface1Method2().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::StaticMethod()._Started.0\) then 
                            \ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::StaticMethod()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::Interface1Method2().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::Interface1Method2().0.runningIndex.0\ := 0;
                            \ComplexTypeHierarchy::StaticMethod().0._Started\ <= true;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::Interface1Method2().0.runningIndex.0\ is 
                            when 0 => 
                                if (\ComplexTypeHierarchy::StaticMethod().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::Interface1Method2().0.runningState.0\ := AfterFinished;
                                    \ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::StaticMethod()._Finished.0\ <= true;
                                    \ComplexTypeHierarchy::StaticMethod().0._Started\ <= false;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::StaticMethod()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::Interface1Method2().0.runningState.0\ := WaitingForStarted;
                            \ComplexTypeHierarchy::Interface1Method2().0.ComplexTypeHierarchy::StaticMethod()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::BaseInterfaceMethod2().0
                case \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::BaseInterfaceMethod2().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\ComplexTypeHierarchy::BaseInterfaceMethod2().0.ComplexTypeHierarchy::StaticMethod()._Started.0\) then 
                            \ComplexTypeHierarchy::BaseInterfaceMethod2().0.ComplexTypeHierarchy::StaticMethod()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::BaseInterfaceMethod2().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::BaseInterfaceMethod2().0.runningIndex.0\ := 0;
                            \ComplexTypeHierarchy::StaticMethod().0._Started\ <= true;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::BaseInterfaceMethod2().0.runningIndex.0\ is 
                            when 0 => 
                                if (\ComplexTypeHierarchy::StaticMethod().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::BaseInterfaceMethod2().0.runningState.0\ := AfterFinished;
                                    \ComplexTypeHierarchy::BaseInterfaceMethod2().0.ComplexTypeHierarchy::StaticMethod()._Finished.0\ <= true;
                                    \ComplexTypeHierarchy::StaticMethod().0._Started\ <= false;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\ComplexTypeHierarchy::BaseInterfaceMethod2().0.ComplexTypeHierarchy::StaticMethod()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::BaseInterfaceMethod2().0.runningState.0\ := WaitingForStarted;
                            \ComplexTypeHierarchy::BaseInterfaceMethod2().0.ComplexTypeHierarchy::StaticMethod()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::PrivateMethod().0
                case \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::PrivateMethod().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\ComplexTypeHierarchy::PrivateMethod().0.ComplexTypeHierarchy::StaticMethod()._Started.0\) then 
                            \ComplexTypeHierarchy::PrivateMethod().0.ComplexTypeHierarchy::StaticMethod()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::PrivateMethod().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::PrivateMethod().0.runningIndex.0\ := 0;
                            \ComplexTypeHierarchy::StaticMethod().0._Started\ <= true;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::PrivateMethod().0.runningIndex.0\ is 
                            when 0 => 
                                if (\ComplexTypeHierarchy::StaticMethod().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::PrivateMethod().0.runningState.0\ := AfterFinished;
                                    \ComplexTypeHierarchy::PrivateMethod().0.ComplexTypeHierarchy::StaticMethod()._Finished.0\ <= true;
                                    \ComplexTypeHierarchy::StaticMethod().0._Started\ <= false;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\ComplexTypeHierarchy::PrivateMethod().0.ComplexTypeHierarchy::StaticMethod()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::StaticMethod().ComplexTypeHierarchy::PrivateMethod().0.runningState.0\ := WaitingForStarted;
                            \ComplexTypeHierarchy::PrivateMethod().0.ComplexTypeHierarchy::StaticMethod()._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::StaticMethod() end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::BaseInterfaceMethod2() start
    \Hast::InternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2()\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2().ComplexTypeHierarchy::Interface2Method1().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2().ComplexTypeHierarchy::Interface2Method1().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2().Hast::ExternalInvocationProxy().runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2().Hast::ExternalInvocationProxy().runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2().ComplexTypeHierarchy::Interface2Method1().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2().ComplexTypeHierarchy::Interface2Method1().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2().Hast::ExternalInvocationProxy().runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2().Hast::ExternalInvocationProxy().runningState.0\ := WaitingForStarted;
                \ComplexTypeHierarchy::Interface2Method1().0.ComplexTypeHierarchy::BaseInterfaceMethod2()._Finished.0\ <= false;
                \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2()._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Interface2Method1().0
                case \Hast::InternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2().ComplexTypeHierarchy::Interface2Method1().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\ComplexTypeHierarchy::Interface2Method1().0.ComplexTypeHierarchy::BaseInterfaceMethod2()._Started.0\) then 
                            \ComplexTypeHierarchy::Interface2Method1().0.ComplexTypeHierarchy::BaseInterfaceMethod2()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2().ComplexTypeHierarchy::Interface2Method1().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2().ComplexTypeHierarchy::Interface2Method1().0.runningIndex.0\ := 0;
                            \ComplexTypeHierarchy::BaseInterfaceMethod2().0._Started\ <= true;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2().ComplexTypeHierarchy::Interface2Method1().0.runningIndex.0\ is 
                            when 0 => 
                                if (\ComplexTypeHierarchy::BaseInterfaceMethod2().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2().ComplexTypeHierarchy::Interface2Method1().0.runningState.0\ := AfterFinished;
                                    \ComplexTypeHierarchy::Interface2Method1().0.ComplexTypeHierarchy::BaseInterfaceMethod2()._Finished.0\ <= true;
                                    \ComplexTypeHierarchy::BaseInterfaceMethod2().0._Started\ <= false;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\ComplexTypeHierarchy::Interface2Method1().0.ComplexTypeHierarchy::BaseInterfaceMethod2()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2().ComplexTypeHierarchy::Interface2Method1().0.runningState.0\ := WaitingForStarted;
                            \ComplexTypeHierarchy::Interface2Method1().0.ComplexTypeHierarchy::BaseInterfaceMethod2()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Void Hast::ExternalInvocationProxy()
                case \Hast::InternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2().Hast::ExternalInvocationProxy().runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Hast::ExternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2()._Started.0\) then 
                            \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2().Hast::ExternalInvocationProxy().runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2().Hast::ExternalInvocationProxy().runningIndex.0\ := 0;
                            \ComplexTypeHierarchy::BaseInterfaceMethod2().0._Started\ <= true;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2().Hast::ExternalInvocationProxy().runningIndex.0\ is 
                            when 0 => 
                                if (\ComplexTypeHierarchy::BaseInterfaceMethod2().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2().Hast::ExternalInvocationProxy().runningState.0\ := AfterFinished;
                                    \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2()._Finished.0\ <= true;
                                    \ComplexTypeHierarchy::BaseInterfaceMethod2().0._Started\ <= false;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Hast::ExternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2().Hast::ExternalInvocationProxy().runningState.0\ := WaitingForStarted;
                            \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::BaseInterfaceMethod2()._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::BaseInterfaceMethod2() end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.StaticClass::StaticMethod() start
    \Hast::InternalInvocationProxy().StaticClass::StaticMethod()\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().StaticClass::StaticMethod().StaticReference::StaticClassUsingMethod().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().StaticClass::StaticMethod().StaticReference::StaticClassUsingMethod().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().StaticClass::StaticMethod().Hast::ExternalInvocationProxy().runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().StaticClass::StaticMethod().Hast::ExternalInvocationProxy().runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().StaticClass::StaticMethod().StaticReference::StaticClassUsingMethod().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().StaticClass::StaticMethod().StaticReference::StaticClassUsingMethod().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().StaticClass::StaticMethod().Hast::ExternalInvocationProxy().runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().StaticClass::StaticMethod().Hast::ExternalInvocationProxy().runningState.0\ := WaitingForStarted;
                \StaticReference::StaticClassUsingMethod().0.StaticClass::StaticMethod()._Finished.0\ <= false;
                \Hast::ExternalInvocationProxy().StaticClass::StaticMethod()._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.Void Hast.TestInputs.ClassStructure2.StaticReference::StaticClassUsingMethod().0
                case \Hast::InternalInvocationProxy().StaticClass::StaticMethod().StaticReference::StaticClassUsingMethod().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\StaticReference::StaticClassUsingMethod().0.StaticClass::StaticMethod()._Started.0\) then 
                            \StaticReference::StaticClassUsingMethod().0.StaticClass::StaticMethod()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().StaticClass::StaticMethod().StaticReference::StaticClassUsingMethod().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().StaticClass::StaticMethod().StaticReference::StaticClassUsingMethod().0.runningIndex.0\ := 0;
                            \StaticClass::StaticMethod().0._Started\ <= true;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().StaticClass::StaticMethod().StaticReference::StaticClassUsingMethod().0.runningIndex.0\ is 
                            when 0 => 
                                if (\StaticClass::StaticMethod().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().StaticClass::StaticMethod().StaticReference::StaticClassUsingMethod().0.runningState.0\ := AfterFinished;
                                    \StaticReference::StaticClassUsingMethod().0.StaticClass::StaticMethod()._Finished.0\ <= true;
                                    \StaticClass::StaticMethod().0._Started\ <= false;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\StaticReference::StaticClassUsingMethod().0.StaticClass::StaticMethod()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().StaticClass::StaticMethod().StaticReference::StaticClassUsingMethod().0.runningState.0\ := WaitingForStarted;
                            \StaticReference::StaticClassUsingMethod().0.StaticClass::StaticMethod()._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Void Hast::ExternalInvocationProxy()
                case \Hast::InternalInvocationProxy().StaticClass::StaticMethod().Hast::ExternalInvocationProxy().runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Hast::ExternalInvocationProxy().StaticClass::StaticMethod()._Started.0\) then 
                            \Hast::ExternalInvocationProxy().StaticClass::StaticMethod()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().StaticClass::StaticMethod().Hast::ExternalInvocationProxy().runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().StaticClass::StaticMethod().Hast::ExternalInvocationProxy().runningIndex.0\ := 0;
                            \StaticClass::StaticMethod().0._Started\ <= true;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().StaticClass::StaticMethod().Hast::ExternalInvocationProxy().runningIndex.0\ is 
                            when 0 => 
                                if (\StaticClass::StaticMethod().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().StaticClass::StaticMethod().Hast::ExternalInvocationProxy().runningState.0\ := AfterFinished;
                                    \Hast::ExternalInvocationProxy().StaticClass::StaticMethod()._Finished.0\ <= true;
                                    \StaticClass::StaticMethod().0._Started\ <= false;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\Hast::ExternalInvocationProxy().StaticClass::StaticMethod()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().StaticClass::StaticMethod().Hast::ExternalInvocationProxy().runningState.0\ := WaitingForStarted;
                            \Hast::ExternalInvocationProxy().StaticClass::StaticMethod()._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.StaticClass::StaticMethod() end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ArrayUsingCases/ArrayHolder::.ctor(System.Int32[]) start
    -- Signal connections for System.Void Hast.TestInputs.Various.ArrayUsingCases::PassArrayToConstructor().0 (#0):
    \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._Started\ <= \ArrayUsingCases::PassArrayToConstructor().0.ArrayUsingCases/ArrayHolder::.ctor(Int32[])._Started.0\;
    \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0.this.parameter.In\ <= \ArrayUsingCases::PassArrayToConstructor().0.ArrayUsingCases/ArrayHolder::.ctor(Int32[]).this.parameter.Out.0\;
    \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0.array.parameter.In\ <= \ArrayUsingCases::PassArrayToConstructor().0.ArrayUsingCases/ArrayHolder::.ctor(Int32[]).array.parameter.Out.0\;
    \ArrayUsingCases::PassArrayToConstructor().0.ArrayUsingCases/ArrayHolder::.ctor(Int32[])._Finished.0\ <= \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0._Finished\;
    \ArrayUsingCases::PassArrayToConstructor().0.ArrayUsingCases/ArrayHolder::.ctor(Int32[]).this.parameter.In.0\ <= \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0.this.parameter.Out\;
    \ArrayUsingCases::PassArrayToConstructor().0.ArrayUsingCases/ArrayHolder::.ctor(Int32[]).array.parameter.In.0\ <= \ArrayUsingCases/ArrayHolder::.ctor(Int32[]).0.array.parameter.Out\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ArrayUsingCases/ArrayHolder::.ctor(System.Int32[]) end


    -- System.Void Hast::InternalInvocationProxy().System.Int32[] Hast.TestInputs.Various.ArrayUsingCases::ArrayProducingMethod(System.Int32) start
    -- Signal connections for System.Void Hast.TestInputs.Various.ArrayUsingCases::PassArrayFromMethod().0 (#0):
    \ArrayUsingCases::ArrayProducingMethod(Int32).0._Started\ <= \ArrayUsingCases::PassArrayFromMethod().0.ArrayUsingCases::ArrayProducingMethod(Int32)._Started.0\;
    \ArrayUsingCases::ArrayProducingMethod(Int32).0.arrayLength.parameter.In\ <= \ArrayUsingCases::PassArrayFromMethod().0.ArrayUsingCases::ArrayProducingMethod(Int32).arrayLength.parameter.Out.0\;
    \ArrayUsingCases::PassArrayFromMethod().0.ArrayUsingCases::ArrayProducingMethod(Int32)._Finished.0\ <= \ArrayUsingCases::ArrayProducingMethod(Int32).0._Finished\;
    \ArrayUsingCases::PassArrayFromMethod().0.ArrayUsingCases::ArrayProducingMethod(Int32).return.0\ <= \ArrayUsingCases::ArrayProducingMethod(Int32).0.return\;
    -- System.Void Hast::InternalInvocationProxy().System.Int32[] Hast.TestInputs.Various.ArrayUsingCases::ArrayProducingMethod(System.Int32) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32[]) start
    \Hast::InternalInvocationProxy().ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).ConstantsUsingCases::ConstantPassingToObject().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).ConstantsUsingCases::ConstantPassingToObject().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                -- Synchronous reset
                \Hast::InternalInvocationProxy().ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).ConstantsUsingCases::ConstantPassingToObject().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).ConstantsUsingCases::ConstantPassingToObject().0.runningState.0\ := WaitingForStarted;
                \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Finished.0\ <= false;
                \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Finished.0\ <= false;
            else 

                -- Invocation handler #0 out of 1 corresponding to System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1).0
                case \Hast::InternalInvocationProxy().ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Started.0\) then 
                            \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.runningIndex.0\ := 0;
                            \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._Started\ <= true;
                            \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.this.parameter.In\ <= \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).this.parameter.Out.0\;
                            \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.array.parameter.In\ <= \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).array.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.runningIndex.0\ is 
                            when 0 => 
                                if (\ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.runningState.0\ := AfterFinished;
                                    \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Finished.0\ <= true;
                                    \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._Started\ <= false;
                                    \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).this.parameter.In.0\ <= \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.this.parameter.Out\;
                                    \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).array.parameter.In.0\ <= \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.array.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.runningState.0\ := WaitingForStarted;
                            \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Finished.0\ <= false;
                        end if;
                end case;


                -- Invocation handler #0 out of 1 corresponding to System.Void Hast.TestInputs.Various.ConstantsUsingCases::ConstantPassingToObject().0
                case \Hast::InternalInvocationProxy().ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).ConstantsUsingCases::ConstantPassingToObject().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Started.0\) then 
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).ConstantsUsingCases::ConstantPassingToObject().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).ConstantsUsingCases::ConstantPassingToObject().0.runningIndex.0\ := 0;
                            \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._Started\ <= true;
                            \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.this.parameter.In\ <= \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).this.parameter.Out.0\;
                            \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.array.parameter.In\ <= \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).array.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).ConstantsUsingCases::ConstantPassingToObject().0.runningIndex.0\ is 
                            when 0 => 
                                if (\ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).ConstantsUsingCases::ConstantPassingToObject().0.runningState.0\ := AfterFinished;
                                    \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Finished.0\ <= true;
                                    \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0._Started\ <= false;
                                    \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).this.parameter.In.0\ <= \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.this.parameter.Out\;
                                    \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).array.parameter.In.0\ <= \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).0.array.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        -- Invoking components need to pull down the Started signal to false.
                        if (\ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[]).ConstantsUsingCases::ConstantPassingToObject().0.runningState.0\ := WaitingForStarted;
                            \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32[])._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32[]) end


    -- System.Void Hast::InternalInvocationProxy().System.Int32 Hast.TestInputs.Various.ConstantsUsingCases::ConstantUsingMethod(System.Int32,System.Int32) start
    -- Signal connections for System.Void Hast.TestInputs.Various.ConstantsUsingCases::ConstantPassingToMethod(System.Int32).0 (#0):
    \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._Started\ <= \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.ConstantsUsingCases::ConstantUsingMethod(Int32,Int32)._Started.0\;
    \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0.input1.parameter.In\ <= \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).input1.parameter.Out.0\;
    \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0.input2.parameter.In\ <= \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).input2.parameter.Out.0\;
    \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.ConstantsUsingCases::ConstantUsingMethod(Int32,Int32)._Finished.0\ <= \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0._Finished\;
    \ConstantsUsingCases::ConstantPassingToMethod(Int32).0.ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).return.0\ <= \ConstantsUsingCases::ConstantUsingMethod(Int32,Int32).0.return\;
    -- System.Void Hast::InternalInvocationProxy().System.Int32 Hast.TestInputs.Various.ConstantsUsingCases::ConstantUsingMethod(System.Int32,System.Int32) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32) start
    -- Signal connections for System.Void Hast.TestInputs.Various.ConstantsUsingCases::ConstantPassingToObject().0 (#0):
    \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._Started\ <= \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32)._Started.0\;
    \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0.this.parameter.In\ <= \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).this.parameter.Out.0\;
    \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0.size.parameter.In\ <= \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).size.parameter.Out.0\;
    \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32)._Finished.0\ <= \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0._Finished\;
    \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).this.parameter.In.0\ <= \ConstantsUsingCases/ArrayHolder1::.ctor(UInt32).0.this.parameter.Out\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(System.UInt32) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1) start
    -- Signal connections for System.Void Hast.TestInputs.Various.ConstantsUsingCases::ConstantPassingToObject().0 (#0):
    \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._Started\ <= \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1)._Started.0\;
    \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.this.parameter.In\ <= \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).this.parameter.Out.0\;
    \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.previous.parameter.In\ <= \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).previous.parameter.Out.0\;
    \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1)._Finished.0\ <= \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0._Finished\;
    \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).this.parameter.In.0\ <= \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.this.parameter.Out\;
    \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).previous.parameter.In.0\ <= \ConstantsUsingCases/ArrayHolder1::.ctor(ConstantsUsingCases/ArrayHolder1).0.previous.parameter.Out\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1::.ctor(Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder1) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder2::.ctor(System.UInt32) start
    -- Signal connections for System.Void Hast.TestInputs.Various.ConstantsUsingCases::ConstantPassingToObject().0 (#0):
    \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._Started\ <= \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32)._Started.0\;
    \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.this.parameter.In\ <= \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).this.parameter.Out.0\;
    \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.size.parameter.In\ <= \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).size.parameter.Out.0\;
    \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32)._Finished.0\ <= \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0._Finished\;
    \ConstantsUsingCases::ConstantPassingToObject().0.ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).this.parameter.In.0\ <= \ConstantsUsingCases/ArrayHolder2::.ctor(UInt32).0.this.parameter.Out\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ConstantsUsingCases/ArrayHolder2::.ctor(System.UInt32) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ObjectUsingCases::VoidMethod(Hast.TestInputs.Various.ObjectUsingCases/MyClass) start
    -- Signal connections for System.Void Hast.TestInputs.Various.ObjectUsingCases::VoidReturn(System.Int32).0 (#0):
    \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._Started\ <= \ObjectUsingCases::VoidReturn(Int32).0.ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass)._Started.0\;
    \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.myClass.parameter.In\ <= \ObjectUsingCases::VoidReturn(Int32).0.ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).myClass.parameter.Out.0\;
    \ObjectUsingCases::VoidReturn(Int32).0.ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass)._Finished.0\ <= \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0._Finished\;
    \ObjectUsingCases::VoidReturn(Int32).0.ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).myClass.parameter.In.0\ <= \ObjectUsingCases::VoidMethod(ObjectUsingCases/MyClass).0.myClass.parameter.Out\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ObjectUsingCases::VoidMethod(Hast.TestInputs.Various.ObjectUsingCases/MyClass) end


    -- System.Void Hast::InternalInvocationProxy().System.Boolean Hast.TestInputs.Various.ParallelCases/Calculator::IsEven() start
    -- Signal connections for System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(System.UInt32).0 (#0):
    \ParallelCases/Calculator::IsEven().0._Started\ <= \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.ParallelCases/Calculator::IsEven()._Started.0\;
    \ParallelCases/Calculator::IsEven().0.this.parameter.In\ <= \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.ParallelCases/Calculator::IsEven().this.parameter.Out.0\;
    \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.ParallelCases/Calculator::IsEven()._Finished.0\ <= \ParallelCases/Calculator::IsEven().0._Finished\;
    \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.ParallelCases/Calculator::IsEven().return.0\ <= \ParallelCases/Calculator::IsEven().0.return\;
    \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.ParallelCases/Calculator::IsEven().this.parameter.In.0\ <= \ParallelCases/Calculator::IsEven().0.this.parameter.Out\;
    -- Signal connections for System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(System.UInt32).1 (#1):
    \ParallelCases/Calculator::IsEven().1._Started\ <= \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.ParallelCases/Calculator::IsEven()._Started.0\;
    \ParallelCases/Calculator::IsEven().1.this.parameter.In\ <= \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.ParallelCases/Calculator::IsEven().this.parameter.Out.0\;
    \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.ParallelCases/Calculator::IsEven()._Finished.0\ <= \ParallelCases/Calculator::IsEven().1._Finished\;
    \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.ParallelCases/Calculator::IsEven().return.0\ <= \ParallelCases/Calculator::IsEven().1.return\;
    \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.ParallelCases/Calculator::IsEven().this.parameter.In.0\ <= \ParallelCases/Calculator::IsEven().1.this.parameter.Out\;
    -- Signal connections for System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(System.UInt32).2 (#2):
    \ParallelCases/Calculator::IsEven().2._Started\ <= \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.ParallelCases/Calculator::IsEven()._Started.0\;
    \ParallelCases/Calculator::IsEven().2.this.parameter.In\ <= \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.ParallelCases/Calculator::IsEven().this.parameter.Out.0\;
    \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.ParallelCases/Calculator::IsEven()._Finished.0\ <= \ParallelCases/Calculator::IsEven().2._Finished\;
    \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.ParallelCases/Calculator::IsEven().return.0\ <= \ParallelCases/Calculator::IsEven().2.return\;
    \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.ParallelCases/Calculator::IsEven().this.parameter.In.0\ <= \ParallelCases/Calculator::IsEven().2.this.parameter.Out\;
    -- System.Void Hast::InternalInvocationProxy().System.Boolean Hast.TestInputs.Various.ParallelCases/Calculator::IsEven() end


    -- System.Void Hast::InternalInvocationProxy().System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(System.UInt32) start
    -- Signal connections for System.Void Hast.TestInputs.Various.ParallelCases::WhenAllWhenAnyAwaitedTasks(System.UInt32).0 (#0):
    \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._Started\ <= \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.0\;
    \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.indexObject.parameter.In\ <= \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).indexObject.parameter.Out.0\;
    \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Finished.0\ <= \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0._Finished\;
    \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).return.0\ <= \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).0.return\;
    -- Signal connections for System.Void Hast.TestInputs.Various.ParallelCases::WhenAllWhenAnyAwaitedTasks(System.UInt32).0 (#1):
    \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._Started\ <= \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.1\;
    \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.indexObject.parameter.In\ <= \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).indexObject.parameter.Out.1\;
    \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Finished.1\ <= \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1._Finished\;
    \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).return.1\ <= \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).1.return\;
    -- Signal connections for System.Void Hast.TestInputs.Various.ParallelCases::WhenAllWhenAnyAwaitedTasks(System.UInt32).0 (#2):
    \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._Started\ <= \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Started.2\;
    \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.indexObject.parameter.In\ <= \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).indexObject.parameter.Out.2\;
    \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32)._Finished.2\ <= \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2._Finished\;
    \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).return.2\ <= \ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(UInt32).2.return\;
    -- System.Void Hast::InternalInvocationProxy().System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass0_0::<WhenAllWhenAnyAwaitedTasks>b__0(System.UInt32) end


    -- System.Void Hast::InternalInvocationProxy().System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(System.UInt32) start
    -- Signal connections for System.Void Hast.TestInputs.Various.ParallelCases::ObjectUsingTasks(System.UInt32).0 (#0):
    \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._Started\ <= \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Started.0\;
    \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.indexObject.parameter.In\ <= \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).indexObject.parameter.Out.0\;
    \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Finished.0\ <= \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0._Finished\;
    \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).return.0\ <= \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).0.return\;
    -- Signal connections for System.Void Hast.TestInputs.Various.ParallelCases::ObjectUsingTasks(System.UInt32).0 (#1):
    \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._Started\ <= \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Started.1\;
    \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.indexObject.parameter.In\ <= \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).indexObject.parameter.Out.1\;
    \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Finished.1\ <= \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1._Finished\;
    \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).return.1\ <= \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).1.return\;
    -- Signal connections for System.Void Hast.TestInputs.Various.ParallelCases::ObjectUsingTasks(System.UInt32).0 (#2):
    \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._Started\ <= \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Started.2\;
    \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.indexObject.parameter.In\ <= \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).indexObject.parameter.Out.2\;
    \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32)._Finished.2\ <= \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2._Finished\;
    \ParallelCases::ObjectUsingTasks(UInt32).0.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).return.2\ <= \ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(UInt32).2.return\;
    -- System.Void Hast::InternalInvocationProxy().System.Boolean Hast.TestInputs.Various.ParallelCases/<>c__DisplayClass1_0::<ObjectUsingTasks>b__0(System.UInt32) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure1.RootClass::VirtualMethod(System.Int32) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \RootClass::VirtualMethod(Int32).0._Started\ <= \Hast::ExternalInvocationProxy().RootClass::VirtualMethod(Int32)._Started.0\;
    \Hast::ExternalInvocationProxy().RootClass::VirtualMethod(Int32)._Finished.0\ <= \RootClass::VirtualMethod(Int32).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure1.RootClass::VirtualMethod(System.Int32) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1() start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._Started\ <= \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1()._Started.0\;
    \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1()._Finished.0\ <= \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1().0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IInterface1.Interface1Method1() end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Interface1Method2() start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \ComplexTypeHierarchy::Interface1Method2().0._Started\ <= \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Interface1Method2()._Started.0\;
    \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Interface1Method2()._Finished.0\ <= \ComplexTypeHierarchy::Interface1Method2().0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Interface1Method2() end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Interface2Method1() start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \ComplexTypeHierarchy::Interface2Method1().0._Started\ <= \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Interface2Method1()._Started.0\;
    \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Interface2Method1()._Finished.0\ <= \ComplexTypeHierarchy::Interface2Method1().0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Interface2Method1() end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1() start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._Started\ <= \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1()._Started.0\;
    \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1()._Finished.0\ <= \ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1().0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::Hast.TestInputs.ClassStructure1.ComplexTypes.IBaseInterface.BaseInterfaceMethod1() end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::NonVirtualNonInterfaceMehod() start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._Started\ <= \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::NonVirtualNonInterfaceMehod()._Started.0\;
    \Hast::ExternalInvocationProxy().ComplexTypeHierarchy::NonVirtualNonInterfaceMehod()._Finished.0\ <= \ComplexTypeHierarchy::NonVirtualNonInterfaceMehod().0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.ComplexTypeHierarchy::NonVirtualNonInterfaceMehod() end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.UnusedDeclarations::UnusedMethod() start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \UnusedDeclarations::UnusedMethod().0._Started\ <= \Hast::ExternalInvocationProxy().UnusedDeclarations::UnusedMethod()._Started.0\;
    \Hast::ExternalInvocationProxy().UnusedDeclarations::UnusedMethod()._Finished.0\ <= \UnusedDeclarations::UnusedMethod().0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure1.ComplexTypes.UnusedDeclarations::UnusedMethod() end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure2.StaticReference::StaticClassUsingMethod() start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \StaticReference::StaticClassUsingMethod().0._Started\ <= \Hast::ExternalInvocationProxy().StaticReference::StaticClassUsingMethod()._Started.0\;
    \Hast::ExternalInvocationProxy().StaticReference::StaticClassUsingMethod()._Finished.0\ <= \StaticReference::StaticClassUsingMethod().0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.ClassStructure2.StaticReference::StaticClassUsingMethod() end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ArrayUsingCases::PassArrayToConstructor() start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \ArrayUsingCases::PassArrayToConstructor().0._Started\ <= \Hast::ExternalInvocationProxy().ArrayUsingCases::PassArrayToConstructor()._Started.0\;
    \Hast::ExternalInvocationProxy().ArrayUsingCases::PassArrayToConstructor()._Finished.0\ <= \ArrayUsingCases::PassArrayToConstructor().0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ArrayUsingCases::PassArrayToConstructor() end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ArrayUsingCases::PassArrayFromMethod() start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \ArrayUsingCases::PassArrayFromMethod().0._Started\ <= \Hast::ExternalInvocationProxy().ArrayUsingCases::PassArrayFromMethod()._Started.0\;
    \Hast::ExternalInvocationProxy().ArrayUsingCases::PassArrayFromMethod()._Finished.0\ <= \ArrayUsingCases::PassArrayFromMethod().0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ArrayUsingCases::PassArrayFromMethod() end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.CastingCases::NumberCasting(System.Int16,System.Int16) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \CastingCases::NumberCasting(Int16,Int16).0._Started\ <= \Hast::ExternalInvocationProxy().CastingCases::NumberCasting(Int16,Int16)._Started.0\;
    \Hast::ExternalInvocationProxy().CastingCases::NumberCasting(Int16,Int16)._Finished.0\ <= \CastingCases::NumberCasting(Int16,Int16).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.CastingCases::NumberCasting(System.Int16,System.Int16) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ConstantsUsingCases::ConstantValuedVariables(System.Int32) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \ConstantsUsingCases::ConstantValuedVariables(Int32).0._Started\ <= \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantValuedVariables(Int32)._Started.0\;
    \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantValuedVariables(Int32)._Finished.0\ <= \ConstantsUsingCases::ConstantValuedVariables(Int32).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ConstantsUsingCases::ConstantValuedVariables(System.Int32) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ConstantsUsingCases::ConstantPassingToMethod(System.Int32) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._Started\ <= \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantPassingToMethod(Int32)._Started.0\;
    \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantPassingToMethod(Int32)._Finished.0\ <= \ConstantsUsingCases::ConstantPassingToMethod(Int32).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ConstantsUsingCases::ConstantPassingToMethod(System.Int32) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ConstantsUsingCases::ConstantPassingToObject() start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \ConstantsUsingCases::ConstantPassingToObject().0._Started\ <= \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantPassingToObject()._Started.0\;
    \Hast::ExternalInvocationProxy().ConstantsUsingCases::ConstantPassingToObject()._Finished.0\ <= \ConstantsUsingCases::ConstantPassingToObject().0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ConstantsUsingCases::ConstantPassingToObject() end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.LoopCases::BreakInLoop(System.Int32) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \LoopCases::BreakInLoop(Int32).0._Started\ <= \Hast::ExternalInvocationProxy().LoopCases::BreakInLoop(Int32)._Started.0\;
    \Hast::ExternalInvocationProxy().LoopCases::BreakInLoop(Int32)._Finished.0\ <= \LoopCases::BreakInLoop(Int32).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.LoopCases::BreakInLoop(System.Int32) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.LoopCases::BreakInLoopInLoop(System.Int32) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \LoopCases::BreakInLoopInLoop(Int32).0._Started\ <= \Hast::ExternalInvocationProxy().LoopCases::BreakInLoopInLoop(Int32)._Started.0\;
    \Hast::ExternalInvocationProxy().LoopCases::BreakInLoopInLoop(Int32)._Finished.0\ <= \LoopCases::BreakInLoopInLoop(Int32).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.LoopCases::BreakInLoopInLoop(System.Int32) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ObjectUsingCases::NullUsage() start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \ObjectUsingCases::NullUsage().0._Started\ <= \Hast::ExternalInvocationProxy().ObjectUsingCases::NullUsage()._Started.0\;
    \Hast::ExternalInvocationProxy().ObjectUsingCases::NullUsage()._Finished.0\ <= \ObjectUsingCases::NullUsage().0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ObjectUsingCases::NullUsage() end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ObjectUsingCases::VoidReturn(System.Int32) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \ObjectUsingCases::VoidReturn(Int32).0._Started\ <= \Hast::ExternalInvocationProxy().ObjectUsingCases::VoidReturn(Int32)._Started.0\;
    \Hast::ExternalInvocationProxy().ObjectUsingCases::VoidReturn(Int32)._Finished.0\ <= \ObjectUsingCases::VoidReturn(Int32).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ObjectUsingCases::VoidReturn(System.Int32) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ParallelCases::WhenAllWhenAnyAwaitedTasks(System.UInt32) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._Started\ <= \Hast::ExternalInvocationProxy().ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32)._Started.0\;
    \Hast::ExternalInvocationProxy().ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32)._Finished.0\ <= \ParallelCases::WhenAllWhenAnyAwaitedTasks(UInt32).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ParallelCases::WhenAllWhenAnyAwaitedTasks(System.UInt32) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ParallelCases::ObjectUsingTasks(System.UInt32) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \ParallelCases::ObjectUsingTasks(UInt32).0._Started\ <= \Hast::ExternalInvocationProxy().ParallelCases::ObjectUsingTasks(UInt32)._Started.0\;
    \Hast::ExternalInvocationProxy().ParallelCases::ObjectUsingTasks(UInt32)._Finished.0\ <= \ParallelCases::ObjectUsingTasks(UInt32).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.ParallelCases::ObjectUsingTasks(System.UInt32) end


    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.UnaryCases::IncrementDecrement(System.Int32) start
    -- Signal connections for System.Void Hast::ExternalInvocationProxy() (#0):
    \UnaryCases::IncrementDecrement(Int32).0._Started\ <= \Hast::ExternalInvocationProxy().UnaryCases::IncrementDecrement(Int32)._Started.0\;
    \Hast::ExternalInvocationProxy().UnaryCases::IncrementDecrement(Int32)._Finished.0\ <= \UnaryCases::IncrementDecrement(Int32).0._Finished\;
    -- System.Void Hast::InternalInvocationProxy().System.Void Hast.TestInputs.Various.UnaryCases::IncrementDecrement(System.Int32) end

end Imp;
