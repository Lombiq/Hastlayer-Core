




library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package TypeConversion is
    function SmartResize(input: unsigned; size: natural) return unsigned;
    function SmartResize(input: signed; size: natural) return signed;
    function ToUnsignedAndExpand(input: signed; size: natural) return unsigned;
end TypeConversion;
        
package body TypeConversion is

    
    
    
    
    
    
    function SmartResize(input: unsigned; size: natural) return unsigned is
    begin
        if (size < input'LENGTH) then
            return input(size - 1 downto 0);
        else
            
            
            
            return resize(input, size);
        end if;
    end SmartResize;

    function SmartResize(input: signed; size: natural) return signed is
    begin
        if (size < input'LENGTH) then
            return input(size - 1 downto 0);
        else
            return resize(input, size);
        end if;
    end SmartResize;

    function ToUnsignedAndExpand(input: signed; size: natural) return unsigned is
        variable result: unsigned(size - 1 downto 0);
    begin
        if (input >= 0) then
            return resize(unsigned(input), size);
        else 
            result := (others => '1');
            result(input'LENGTH - 1 downto 0) := unsigned(input);
            return result;
        end if;
    end ToUnsignedAndExpand;

end TypeConversion;


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
        
package SimpleMemory is
    
    function ConvertUInt32ToStdLogicVector(input: unsigned(31 downto 0)) return std_logic_vector;
    function ConvertStdLogicVectorToUInt32(input : std_logic_vector) return unsigned;
        
    function ConvertBooleanToStdLogicVector(input: boolean) return std_logic_vector;
    function ConvertStdLogicVectorToBoolean(input : std_logic_vector) return boolean;
        
    function ConvertInt32ToStdLogicVector(input: signed(31 downto 0)) return std_logic_vector;
    function ConvertStdLogicVectorToInt32(input : std_logic_vector) return signed;
end SimpleMemory;
        
package body SimpleMemory is

    function ConvertUInt32ToStdLogicVector(input: unsigned(31 downto 0)) return std_logic_vector is
    begin
        return std_logic_vector(input);
    end ConvertUInt32ToStdLogicVector;
    
    function ConvertStdLogicVectorToUInt32(input : std_logic_vector) return unsigned is
    begin
        return unsigned(input);
    end ConvertStdLogicVectorToUInt32;
    
    function ConvertBooleanToStdLogicVector(input: boolean) return std_logic_vector is 
    begin
        case input is
            when true => return X"FFFFFFFF";
            when false => return X"00000000";
            when others => return X"00000000";
        end case;
    end ConvertBooleanToStdLogicVector;

    function ConvertStdLogicVectorToBoolean(input : std_logic_vector) return boolean is 
    begin
        
        return not(input = X"00000000");
    end ConvertStdLogicVectorToBoolean;

    function ConvertInt32ToStdLogicVector(input: signed(31 downto 0)) return std_logic_vector is
    begin
        return std_logic_vector(input);
    end ConvertInt32ToStdLogicVector;

    function ConvertStdLogicVectorToInt32(input : std_logic_vector) return signed is
    begin
        return signed(input);
    end ConvertStdLogicVectorToInt32;

end SimpleMemory;


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.TypeConversion.all;
library work;
use work.SimpleMemory.all;

entity Hast_IP is 
    port(
        \DataIn\: In std_logic_vector(31 downto 0);
        \DataOut\: Out std_logic_vector(31 downto 0);
        \CellIndex\: Out integer;
        \ReadEnable\: Out boolean;
        \WriteEnable\: Out boolean;
        \ReadsDone\: In boolean;
        \WritesDone\: In boolean;
        \MemberId\: In integer;
        \Reset\: In std_logic;
        \Started\: In boolean;
        \Finished\: Out boolean;
        \Clock\: In std_logic
    );
    
    
    

    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    

end Hast_IP;

architecture Imp of Hast_IP is 
    
    
    
    
    
    
    
    
    

    
    attribute altera_attribute: string;
    attribute altera_attribute of Imp: architecture is "-name SDC_STATEMENT ""set_multicycle_path 8 -setup -to {*Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._StateMachine:Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.0[*]}"";-name SDC_STATEMENT ""set_multicycle_path 7 -hold -to {*Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._StateMachine:Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.0[*]}"";-name SDC_STATEMENT ""set_multicycle_path 8 -setup -to {*Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._StateMachine:Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.1[*]}"";-name SDC_STATEMENT ""set_multicycle_path 7 -hold -to {*Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._StateMachine:Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.1[*]}""";


    
    type \Lombiq.Arithmetics.Posit32\ is record 
        \IsNull\: boolean;
        \PositBits\: unsigned(31 downto 0);
    end record;
    type \Lombiq.Arithmetics.Posit32_Array\ is array (integer range <>) of \Lombiq.Arithmetics.Posit32\;
    type \unsigned64_Array\ is array (integer range <>) of unsigned(63 downto 0);
    type \Lombiq.Arithmetics.Quire\ is record 
        \IsNull\: boolean;
        \Size\: unsigned(15 downto 0);
        \SegmentCount\: unsigned(15 downto 0);
        \Segments\: \unsigned64_Array\(0 to 7);
    end record;
    


    
    
    type \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._States\ is (
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_0\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_1\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_2\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_3\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_4\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_5\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_6\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_7\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_8\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_9\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_10\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_11\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_12\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_13\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_14\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_15\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_16\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_17\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_18\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_19\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_20\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_21\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_22\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_23\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_24\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_25\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_26\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_27\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_28\);
    
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._Finished\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.DataOut\: std_logic_vector(31 downto 0) := (others => '0');
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.ReadEnable\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.WriteEnable\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).this.parameter.Out.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).value.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Started.0\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32).x.parameter.Out.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Started.0\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).this.parameter.Out.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).bits.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).fromBitMask.parameter.Out.0\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean)._Started.0\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).posits.parameter.Out.0\: \Lombiq.Arithmetics.Posit32_Array\(0 to 159);
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).startingValue.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire)._Started.0\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).this.parameter.Out.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).q.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire)._Started.0\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._Started\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).this.parameter.In.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Finished.0\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32).return.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).this.parameter.In.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean)._Finished.0\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).posits.parameter.In.0\: \Lombiq.Arithmetics.Posit32_Array\(0 to 159);
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).startingValue.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire)._Finished.0\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).return.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).this.parameter.In.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).q.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire)._Finished.0\: boolean := false;
    


    
    
    type \Posit32::.ctor(UInt32,Boolean).0._States\ is (
        \Posit32::.ctor(UInt32,Boolean).0._State_0\, 
        \Posit32::.ctor(UInt32,Boolean).0._State_1\, 
        \Posit32::.ctor(UInt32,Boolean).0._State_2\);
    
    Signal \Posit32::.ctor(UInt32,Boolean).0._Finished\: boolean := false;
    Signal \Posit32::.ctor(UInt32,Boolean).0.this.parameter.Out\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::.ctor(UInt32,Boolean).0._Started\: boolean := false;
    Signal \Posit32::.ctor(UInt32,Boolean).0.this.parameter.In\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::.ctor(UInt32,Boolean).0.bits.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::.ctor(UInt32,Boolean).0.fromBitMask.parameter.In\: boolean := false;
    


    
    
    type \Posit32::.ctor(Quire).0._States\ is (
        \Posit32::.ctor(Quire).0._State_0\, 
        \Posit32::.ctor(Quire).0._State_1\, 
        \Posit32::.ctor(Quire).0._State_2\, 
        \Posit32::.ctor(Quire).0._State_3\, 
        \Posit32::.ctor(Quire).0._State_4\, 
        \Posit32::.ctor(Quire).0._State_5\, 
        \Posit32::.ctor(Quire).0._State_6\, 
        \Posit32::.ctor(Quire).0._State_7\, 
        \Posit32::.ctor(Quire).0._State_8\, 
        \Posit32::.ctor(Quire).0._State_9\, 
        \Posit32::.ctor(Quire).0._State_10\, 
        \Posit32::.ctor(Quire).0._State_11\, 
        \Posit32::.ctor(Quire).0._State_12\, 
        \Posit32::.ctor(Quire).0._State_13\, 
        \Posit32::.ctor(Quire).0._State_14\, 
        \Posit32::.ctor(Quire).0._State_15\, 
        \Posit32::.ctor(Quire).0._State_16\, 
        \Posit32::.ctor(Quire).0._State_17\, 
        \Posit32::.ctor(Quire).0._State_18\, 
        \Posit32::.ctor(Quire).0._State_19\, 
        \Posit32::.ctor(Quire).0._State_20\, 
        \Posit32::.ctor(Quire).0._State_21\, 
        \Posit32::.ctor(Quire).0._State_22\, 
        \Posit32::.ctor(Quire).0._State_23\, 
        \Posit32::.ctor(Quire).0._State_24\);
    
    Signal \Posit32::.ctor(Quire).0._Finished\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.this.parameter.Out\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::.ctor(Quire).0.q.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).right.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).x.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire).q.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire)._Started.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).left.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).right.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32)._Started.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire).x.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire)._Started.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).signBit.parameter.Out.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).regimeKValue.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).exponentBits.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).fractionBits.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32)._Started.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0._Started\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.this.parameter.In\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::.ctor(Quire).0.q.parameter.In\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Finished.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).return.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).x.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Finished.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).return.0\: unsigned(63 downto 0) := to_unsigned(0, 64);
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire).q.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire)._Finished.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire).return.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).left.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32)._Finished.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).return.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).return.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire).x.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire)._Finished.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32)._Finished.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    


    
    
    type \Posit32::.ctor(UInt32).0._States\ is (
        \Posit32::.ctor(UInt32).0._State_0\, 
        \Posit32::.ctor(UInt32).0._State_1\, 
        \Posit32::.ctor(UInt32).0._State_2\);
    
    Signal \Posit32::.ctor(UInt32).0._Finished\: boolean := false;
    Signal \Posit32::.ctor(UInt32).0.this.parameter.Out\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::.ctor(UInt32).0._Started\: boolean := false;
    Signal \Posit32::.ctor(UInt32).0.this.parameter.In\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::.ctor(UInt32).0.value.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    


    
    
    type \Posit32::.ctor(Int32).0._States\ is (
        \Posit32::.ctor(Int32).0._State_0\, 
        \Posit32::.ctor(Int32).0._State_1\, 
        \Posit32::.ctor(Int32).0._State_2\, 
        \Posit32::.ctor(Int32).0._State_3\);
    
    Signal \Posit32::.ctor(Int32).0._Finished\: boolean := false;
    Signal \Posit32::.ctor(Int32).0.this.parameter.Out\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32).this.parameter.Out.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32).value.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32)._Started.0\: boolean := false;
    Signal \Posit32::.ctor(Int32).0._Started\: boolean := false;
    Signal \Posit32::.ctor(Int32).0.this.parameter.In\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::.ctor(Int32).0.value.parameter.In\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32).this.parameter.In.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32)._Finished.0\: boolean := false;
    


    
    
    type \Posit32::IsNaN().0._States\ is (
        \Posit32::IsNaN().0._State_0\, 
        \Posit32::IsNaN().0._State_1\, 
        \Posit32::IsNaN().0._State_2\);
    
    Signal \Posit32::IsNaN().0._Finished\: boolean := false;
    Signal \Posit32::IsNaN().0.return\: boolean := false;
    Signal \Posit32::IsNaN().0._Started\: boolean := false;
    Signal \Posit32::IsNaN().0.this.parameter.In\: \Lombiq.Arithmetics.Posit32\;
    


    
    
    type \Posit32::EncodeRegimeBits(Int32).0._States\ is (
        \Posit32::EncodeRegimeBits(Int32).0._State_0\, 
        \Posit32::EncodeRegimeBits(Int32).0._State_1\, 
        \Posit32::EncodeRegimeBits(Int32).0._State_2\, 
        \Posit32::EncodeRegimeBits(Int32).0._State_3\, 
        \Posit32::EncodeRegimeBits(Int32).0._State_4\, 
        \Posit32::EncodeRegimeBits(Int32).0._State_5\, 
        \Posit32::EncodeRegimeBits(Int32).0._State_6\, 
        \Posit32::EncodeRegimeBits(Int32).0._State_7\);
    
    Signal \Posit32::EncodeRegimeBits(Int32).0._Finished\: boolean := false;
    Signal \Posit32::EncodeRegimeBits(Int32).0.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::EncodeRegimeBits(Int32).0.Posit32::GetMostSignificantOnePosition(UInt32).bits.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::EncodeRegimeBits(Int32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Started.0\: boolean := false;
    Signal \Posit32::EncodeRegimeBits(Int32).0._Started\: boolean := false;
    Signal \Posit32::EncodeRegimeBits(Int32).0.regimeKValue.parameter.In\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Posit32::EncodeRegimeBits(Int32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Finished.0\: boolean := false;
    Signal \Posit32::EncodeRegimeBits(Int32).0.Posit32::GetMostSignificantOnePosition(UInt32).return.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
    


    
    
    type \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._States\ is (
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_0\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_1\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_2\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_3\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_4\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_5\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_6\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_7\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_8\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_9\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_10\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_11\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_12\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_13\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_14\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_15\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_16\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_17\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_18\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_19\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_20\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_21\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_22\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_23\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_24\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_25\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_26\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_27\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_28\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_29\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_30\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_31\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_32\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_33\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_34\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_35\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_36\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_37\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_38\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_39\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_40\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_41\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_42\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_43\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_44\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_45\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_46\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_47\);
    
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._Finished\: boolean := false;
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::EncodeRegimeBits(Int32).regimeKValue.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::EncodeRegimeBits(Int32)._Started.0\: boolean := false;
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte).bits.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte).startingPosition.parameter.Out.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\: boolean := false;
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32).bits.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32)._Started.0\: boolean := false;
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetMostSignificantOnePosition(UInt32).bits.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Started.0\: boolean := false;
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::SetZero(UInt32,UInt16).bits.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::SetZero(UInt32,UInt16).index.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::SetZero(UInt32,UInt16)._Started.0\: boolean := false;
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._Started\: boolean := false;
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.signBit.parameter.In\: boolean := false;
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.regimeKValue.parameter.In\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::EncodeRegimeBits(Int32)._Finished.0\: boolean := false;
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::EncodeRegimeBits(Int32).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\: boolean := false;
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte).return.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32)._Finished.0\: boolean := false;
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Finished.0\: boolean := false;
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetMostSignificantOnePosition(UInt32).return.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::SetZero(UInt32,UInt16)._Finished.0\: boolean := false;
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::SetZero(UInt32,UInt16).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    


    
    
    type \Posit32::GetRegimeKValue().0._States\ is (
        \Posit32::GetRegimeKValue().0._State_0\, 
        \Posit32::GetRegimeKValue().0._State_1\, 
        \Posit32::GetRegimeKValue().0._State_2\, 
        \Posit32::GetRegimeKValue().0._State_3\);
    
    Signal \Posit32::GetRegimeKValue().0._Finished\: boolean := false;
    Signal \Posit32::GetRegimeKValue().0.return\: signed(7 downto 0) := to_signed(0, 8);
    Signal \Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte).bits.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte).startingPosition.parameter.Out.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
    Signal \Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\: boolean := false;
    Signal \Posit32::GetRegimeKValue().0._Started\: boolean := false;
    Signal \Posit32::GetRegimeKValue().0.this.parameter.In\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\: boolean := false;
    Signal \Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte).return.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
    


    
    
    type \Posit32::CalculateScaleFactor().0._States\ is (
        \Posit32::CalculateScaleFactor().0._State_0\, 
        \Posit32::CalculateScaleFactor().0._State_1\, 
        \Posit32::CalculateScaleFactor().0._State_2\, 
        \Posit32::CalculateScaleFactor().0._State_3\, 
        \Posit32::CalculateScaleFactor().0._State_4\, 
        \Posit32::CalculateScaleFactor().0._State_5\, 
        \Posit32::CalculateScaleFactor().0._State_6\, 
        \Posit32::CalculateScaleFactor().0._State_7\);
    
    Signal \Posit32::CalculateScaleFactor().0._Finished\: boolean := false;
    Signal \Posit32::CalculateScaleFactor().0.return\: signed(15 downto 0) := to_signed(0, 16);
    Signal \Posit32::CalculateScaleFactor().0.Posit32::GetRegimeKValue().this.parameter.Out.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::CalculateScaleFactor().0.Posit32::GetRegimeKValue()._Started.0\: boolean := false;
    Signal \Posit32::CalculateScaleFactor().0.Posit32::GetExponentValue().this.parameter.Out.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::CalculateScaleFactor().0.Posit32::GetExponentValue()._Started.0\: boolean := false;
    Signal \Posit32::CalculateScaleFactor().0._Started\: boolean := false;
    Signal \Posit32::CalculateScaleFactor().0.this.parameter.In\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::CalculateScaleFactor().0.Posit32::GetRegimeKValue()._Finished.0\: boolean := false;
    Signal \Posit32::CalculateScaleFactor().0.Posit32::GetRegimeKValue().return.0\: signed(7 downto 0) := to_signed(0, 8);
    Signal \Posit32::CalculateScaleFactor().0.Posit32::GetExponentValue()._Finished.0\: boolean := false;
    Signal \Posit32::CalculateScaleFactor().0.Posit32::GetExponentValue().return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    


    
    
    type \Posit32::ExponentSize().0._States\ is (
        \Posit32::ExponentSize().0._State_0\, 
        \Posit32::ExponentSize().0._State_1\, 
        \Posit32::ExponentSize().0._State_2\, 
        \Posit32::ExponentSize().0._State_3\, 
        \Posit32::ExponentSize().0._State_4\, 
        \Posit32::ExponentSize().0._State_5\, 
        \Posit32::ExponentSize().0._State_6\, 
        \Posit32::ExponentSize().0._State_7\, 
        \Posit32::ExponentSize().0._State_8\, 
        \Posit32::ExponentSize().0._State_9\);
    
    Signal \Posit32::ExponentSize().0._Finished\: boolean := false;
    Signal \Posit32::ExponentSize().0.return\: unsigned(7 downto 0) := to_unsigned(0, 8);
    Signal \Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte).bits.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte).startingPosition.parameter.Out.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
    Signal \Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\: boolean := false;
    Signal \Posit32::ExponentSize().0._Started\: boolean := false;
    Signal \Posit32::ExponentSize().0.this.parameter.In\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\: boolean := false;
    Signal \Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte).return.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
    


    
    
    type \Posit32::GetExponentValue().0._States\ is (
        \Posit32::GetExponentValue().0._State_0\, 
        \Posit32::GetExponentValue().0._State_1\, 
        \Posit32::GetExponentValue().0._State_2\, 
        \Posit32::GetExponentValue().0._State_3\, 
        \Posit32::GetExponentValue().0._State_4\, 
        \Posit32::GetExponentValue().0._State_5\, 
        \Posit32::GetExponentValue().0._State_6\, 
        \Posit32::GetExponentValue().0._State_7\, 
        \Posit32::GetExponentValue().0._State_8\, 
        \Posit32::GetExponentValue().0._State_9\);
    
    Signal \Posit32::GetExponentValue().0._Finished\: boolean := false;
    Signal \Posit32::GetExponentValue().0.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::GetExponentValue().0.Posit32::ExponentSize().this.parameter.Out.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::GetExponentValue().0.Posit32::ExponentSize()._Started.0\: boolean := false;
    Signal \Posit32::GetExponentValue().0.Posit32::FractionSize().this.parameter.Out.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::GetExponentValue().0.Posit32::FractionSize()._Started.0\: boolean := false;
    Signal \Posit32::GetExponentValue().0._Started\: boolean := false;
    Signal \Posit32::GetExponentValue().0.this.parameter.In\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::GetExponentValue().0.Posit32::ExponentSize()._Finished.0\: boolean := false;
    Signal \Posit32::GetExponentValue().0.Posit32::ExponentSize().return.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
    Signal \Posit32::GetExponentValue().0.Posit32::FractionSize()._Finished.0\: boolean := false;
    Signal \Posit32::GetExponentValue().0.Posit32::FractionSize().return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    


    
    
    type \Posit32::FractionSize().0._States\ is (
        \Posit32::FractionSize().0._State_0\, 
        \Posit32::FractionSize().0._State_1\, 
        \Posit32::FractionSize().0._State_2\, 
        \Posit32::FractionSize().0._State_3\, 
        \Posit32::FractionSize().0._State_4\, 
        \Posit32::FractionSize().0._State_5\, 
        \Posit32::FractionSize().0._State_6\, 
        \Posit32::FractionSize().0._State_7\);
    
    Signal \Posit32::FractionSize().0._Finished\: boolean := false;
    Signal \Posit32::FractionSize().0.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte).bits.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte).startingPosition.parameter.Out.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
    Signal \Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\: boolean := false;
    Signal \Posit32::FractionSize().0._Started\: boolean := false;
    Signal \Posit32::FractionSize().0.this.parameter.In\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\: boolean := false;
    Signal \Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte).return.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
    


    
    
    type \Posit32::FractionWithHiddenBit().0._States\ is (
        \Posit32::FractionWithHiddenBit().0._State_0\, 
        \Posit32::FractionWithHiddenBit().0._State_1\, 
        \Posit32::FractionWithHiddenBit().0._State_2\, 
        \Posit32::FractionWithHiddenBit().0._State_3\, 
        \Posit32::FractionWithHiddenBit().0._State_4\, 
        \Posit32::FractionWithHiddenBit().0._State_5\, 
        \Posit32::FractionWithHiddenBit().0._State_6\, 
        \Posit32::FractionWithHiddenBit().0._State_7\, 
        \Posit32::FractionWithHiddenBit().0._State_8\, 
        \Posit32::FractionWithHiddenBit().0._State_9\, 
        \Posit32::FractionWithHiddenBit().0._State_10\);
    
    Signal \Posit32::FractionWithHiddenBit().0._Finished\: boolean := false;
    Signal \Posit32::FractionWithHiddenBit().0.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::FractionWithHiddenBit().0.Posit32::FractionSize().this.parameter.Out.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::FractionWithHiddenBit().0.Posit32::FractionSize()._Started.0\: boolean := false;
    Signal \Posit32::FractionWithHiddenBit().0.Posit32::SetOne(UInt32,UInt16).this.parameter.Out.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::FractionWithHiddenBit().0.Posit32::SetOne(UInt32,UInt16).bits.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::FractionWithHiddenBit().0.Posit32::SetOne(UInt32,UInt16).index.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Posit32::FractionWithHiddenBit().0.Posit32::SetOne(UInt32,UInt16)._Started.0\: boolean := false;
    Signal \Posit32::FractionWithHiddenBit().0._Started\: boolean := false;
    Signal \Posit32::FractionWithHiddenBit().0.this.parameter.In\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::FractionWithHiddenBit().0.Posit32::FractionSize()._Finished.0\: boolean := false;
    Signal \Posit32::FractionWithHiddenBit().0.Posit32::FractionSize().return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::FractionWithHiddenBit().0.Posit32::SetOne(UInt32,UInt16)._Finished.0\: boolean := false;
    Signal \Posit32::FractionWithHiddenBit().0.Posit32::SetOne(UInt32,UInt16).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    


    
    
    type \Posit32::GetMostSignificantOnePosition(UInt32).0._States\ is (
        \Posit32::GetMostSignificantOnePosition(UInt32).0._State_0\, 
        \Posit32::GetMostSignificantOnePosition(UInt32).0._State_1\, 
        \Posit32::GetMostSignificantOnePosition(UInt32).0._State_2\, 
        \Posit32::GetMostSignificantOnePosition(UInt32).0._State_3\, 
        \Posit32::GetMostSignificantOnePosition(UInt32).0._State_4\, 
        \Posit32::GetMostSignificantOnePosition(UInt32).0._State_5\);
    
    Signal \Posit32::GetMostSignificantOnePosition(UInt32).0._Finished\: boolean := false;
    Signal \Posit32::GetMostSignificantOnePosition(UInt32).0.return\: unsigned(7 downto 0) := to_unsigned(0, 8);
    Signal \Posit32::GetMostSignificantOnePosition(UInt32).0._Started\: boolean := false;
    Signal \Posit32::GetMostSignificantOnePosition(UInt32).0.bits.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    


    
    
    type \Posit32::SetOne(UInt32,UInt16).0._States\ is (
        \Posit32::SetOne(UInt32,UInt16).0._State_0\, 
        \Posit32::SetOne(UInt32,UInt16).0._State_1\, 
        \Posit32::SetOne(UInt32,UInt16).0._State_2\);
    
    Signal \Posit32::SetOne(UInt32,UInt16).0._Finished\: boolean := false;
    Signal \Posit32::SetOne(UInt32,UInt16).0.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::SetOne(UInt32,UInt16).0._Started\: boolean := false;
    Signal \Posit32::SetOne(UInt32,UInt16).0.this.parameter.In\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::SetOne(UInt32,UInt16).0.bits.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::SetOne(UInt32,UInt16).0.index.parameter.In\: unsigned(15 downto 0) := to_unsigned(0, 16);
    


    
    
    type \Posit32::SetZero(UInt32,UInt16).0._States\ is (
        \Posit32::SetZero(UInt32,UInt16).0._State_0\, 
        \Posit32::SetZero(UInt32,UInt16).0._State_1\, 
        \Posit32::SetZero(UInt32,UInt16).0._State_2\);
    
    Signal \Posit32::SetZero(UInt32,UInt16).0._Finished\: boolean := false;
    Signal \Posit32::SetZero(UInt32,UInt16).0.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::SetZero(UInt32,UInt16).0._Started\: boolean := false;
    Signal \Posit32::SetZero(UInt32,UInt16).0.bits.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::SetZero(UInt32,UInt16).0.index.parameter.In\: unsigned(15 downto 0) := to_unsigned(0, 16);
    


    
    
    type \Posit32::LengthOfRunOfBits(UInt32,Byte).0._States\ is (
        \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_0\, 
        \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_1\, 
        \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_2\, 
        \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_3\, 
        \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_4\, 
        \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_5\, 
        \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_6\);
    
    Signal \Posit32::LengthOfRunOfBits(UInt32,Byte).0._Finished\: boolean := false;
    Signal \Posit32::LengthOfRunOfBits(UInt32,Byte).0.return\: unsigned(7 downto 0) := to_unsigned(0, 8);
    Signal \Posit32::LengthOfRunOfBits(UInt32,Byte).0._Started\: boolean := false;
    Signal \Posit32::LengthOfRunOfBits(UInt32,Byte).0.bits.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::LengthOfRunOfBits(UInt32,Byte).0.startingPosition.parameter.In\: unsigned(7 downto 0) := to_unsigned(0, 8);
    


    
    
    type \Posit32::GetTwosComplement(UInt32).0._States\ is (
        \Posit32::GetTwosComplement(UInt32).0._State_0\, 
        \Posit32::GetTwosComplement(UInt32).0._State_1\, 
        \Posit32::GetTwosComplement(UInt32).0._State_2\);
    
    Signal \Posit32::GetTwosComplement(UInt32).0._Finished\: boolean := false;
    Signal \Posit32::GetTwosComplement(UInt32).0.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::GetTwosComplement(UInt32).0._Started\: boolean := false;
    Signal \Posit32::GetTwosComplement(UInt32).0.bits.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    


    
    
    type \Posit32::FusedSum(Posit32[],Quire).0._States\ is (
        \Posit32::FusedSum(Posit32[],Quire).0._State_0\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_1\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_2\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_3\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_4\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_5\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_6\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_7\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_8\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_9\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_10\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_11\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_12\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_13\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_14\);
    
    Signal \Posit32::FusedSum(Posit32[],Quire).0._Finished\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.return\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.posits.parameter.Out\: \Lombiq.Arithmetics.Posit32_Array\(0 to 159);
    Signal \Posit32::FusedSum(Posit32[],Quire).0.startingValue.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).this.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).firstSegment.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Started.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).left.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).right.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire)._Started.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Posit32::IsNaN().this.parameter.Out.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Posit32::IsNaN()._Started.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32).x.parameter.Out.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Started.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0._Started\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.posits.parameter.In\: \Lombiq.Arithmetics.Posit32_Array\(0 to 159);
    Signal \Posit32::FusedSum(Posit32[],Quire).0.startingValue.parameter.In\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).this.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Finished.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).return.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).left.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).right.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire)._Finished.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).return.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Posit32::IsNaN()._Finished.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Posit32::IsNaN().return.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32).return.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).return.0\: \Lombiq.Arithmetics.Quire\;
    


    
    
    type \Quire Posit32::op_Explicit(Posit32).0._States\ is (
        \Quire Posit32::op_Explicit(Posit32).0._State_0\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_1\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_2\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_3\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_4\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_5\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_6\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_7\);
    
    Signal \Quire Posit32::op_Explicit(Posit32).0._Finished\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0.return\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionWithHiddenBit().this.parameter.Out.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionWithHiddenBit()._Started.0\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionSize().this.parameter.Out.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionSize()._Started.0\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Posit32::CalculateScaleFactor().this.parameter.Out.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Posit32::CalculateScaleFactor()._Started.0\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0._Started\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0.x.parameter.In\: \Lombiq.Arithmetics.Posit32\;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionWithHiddenBit()._Finished.0\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionWithHiddenBit().return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionSize()._Finished.0\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionSize().return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Quire Posit32::op_Explicit(Posit32).0.Posit32::CalculateScaleFactor()._Finished.0\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Posit32::CalculateScaleFactor().return.0\: signed(15 downto 0) := to_signed(0, 16);
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).return.0\: \Lombiq.Arithmetics.Quire\;
    


    
    
    type \Quire::.ctor(UInt64[],UInt16).0._States\ is (
        \Quire::.ctor(UInt64[],UInt16).0._State_0\, 
        \Quire::.ctor(UInt64[],UInt16).0._State_1\, 
        \Quire::.ctor(UInt64[],UInt16).0._State_2\, 
        \Quire::.ctor(UInt64[],UInt16).0._State_3\, 
        \Quire::.ctor(UInt64[],UInt16).0._State_4\);
    
    Signal \Quire::.ctor(UInt64[],UInt16).0._Finished\: boolean := false;
    Signal \Quire::.ctor(UInt64[],UInt16).0.this.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.Out\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
    Signal \Quire::.ctor(UInt64[],UInt16).0._Started\: boolean := false;
    Signal \Quire::.ctor(UInt64[],UInt16).0.this.parameter.In\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.In\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
    Signal \Quire::.ctor(UInt64[],UInt16).0.size.parameter.In\: unsigned(15 downto 0) := to_unsigned(0, 16);
    


    
    
    type \Quire::.ctor(UInt32,UInt16).0._States\ is (
        \Quire::.ctor(UInt32,UInt16).0._State_0\, 
        \Quire::.ctor(UInt32,UInt16).0._State_1\, 
        \Quire::.ctor(UInt32,UInt16).0._State_2\, 
        \Quire::.ctor(UInt32,UInt16).0._State_3\, 
        \Quire::.ctor(UInt32,UInt16).0._State_4\, 
        \Quire::.ctor(UInt32,UInt16).0._State_5\, 
        \Quire::.ctor(UInt32,UInt16).0._State_6\, 
        \Quire::.ctor(UInt32,UInt16).0._State_7\, 
        \Quire::.ctor(UInt32,UInt16).0._State_8\);
    
    Signal \Quire::.ctor(UInt32,UInt16).0._Finished\: boolean := false;
    Signal \Quire::.ctor(UInt32,UInt16).0.this.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire::.ctor(UInt32,UInt16).0._Started\: boolean := false;
    Signal \Quire::.ctor(UInt32,UInt16).0.this.parameter.In\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire::.ctor(UInt32,UInt16).0.firstSegment.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Quire::.ctor(UInt32,UInt16).0.size.parameter.In\: unsigned(15 downto 0) := to_unsigned(0, 16);
    


    
    
    type \Quire Quire::op_Addition(Quire,Quire).0._States\ is (
        \Quire Quire::op_Addition(Quire,Quire).0._State_0\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_1\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_2\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_3\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_4\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_5\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_6\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_7\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_8\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_9\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_10\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_11\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_12\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_13\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_14\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_15\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_16\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_17\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_18\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_19\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_20\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_21\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_22\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_23\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_24\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_25\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_26\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_27\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_28\);
    
    Signal \Quire Quire::op_Addition(Quire,Quire).0._Finished\: boolean := false;
    Signal \Quire Quire::op_Addition(Quire,Quire).0.return\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,Quire).0.left.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,Quire).0.right.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
    Signal \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Started.0\: boolean := false;
    Signal \Quire Quire::op_Addition(Quire,Quire).0._Started\: boolean := false;
    Signal \Quire Quire::op_Addition(Quire,Quire).0.left.parameter.In\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,Quire).0.right.parameter.In\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
    Signal \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\: boolean := false;
    


    
    
    type \Quire Quire::op_Addition(Quire,UInt32).0._States\ is (
        \Quire Quire::op_Addition(Quire,UInt32).0._State_0\, 
        \Quire Quire::op_Addition(Quire,UInt32).0._State_1\, 
        \Quire Quire::op_Addition(Quire,UInt32).0._State_2\, 
        \Quire Quire::op_Addition(Quire,UInt32).0._State_3\, 
        \Quire Quire::op_Addition(Quire,UInt32).0._State_4\);
    
    Signal \Quire Quire::op_Addition(Quire,UInt32).0._Finished\: boolean := false;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.return\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.left.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).this.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).firstSegment.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Started.0\: boolean := false;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\: boolean := false;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0._Started\: boolean := false;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.left.parameter.In\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.right.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).this.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Finished.0\: boolean := false;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\: boolean := false;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).return.0\: \Lombiq.Arithmetics.Quire\;
    


    
    
    type \Quire Quire::op_OnesComplement(Quire).0._States\ is (
        \Quire Quire::op_OnesComplement(Quire).0._State_0\, 
        \Quire Quire::op_OnesComplement(Quire).0._State_1\, 
        \Quire Quire::op_OnesComplement(Quire).0._State_2\, 
        \Quire Quire::op_OnesComplement(Quire).0._State_3\, 
        \Quire Quire::op_OnesComplement(Quire).0._State_4\, 
        \Quire Quire::op_OnesComplement(Quire).0._State_5\);
    
    Signal \Quire Quire::op_OnesComplement(Quire).0._Finished\: boolean := false;
    Signal \Quire Quire::op_OnesComplement(Quire).0.return\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_OnesComplement(Quire).0.q.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_OnesComplement(Quire).0._Started\: boolean := false;
    Signal \Quire Quire::op_OnesComplement(Quire).0.q.parameter.In\: \Lombiq.Arithmetics.Quire\;
    


    
    
    type \Boolean Quire::op_Equality(Quire,Quire).0._States\ is (
        \Boolean Quire::op_Equality(Quire,Quire).0._State_0\, 
        \Boolean Quire::op_Equality(Quire,Quire).0._State_1\, 
        \Boolean Quire::op_Equality(Quire,Quire).0._State_2\, 
        \Boolean Quire::op_Equality(Quire,Quire).0._State_3\, 
        \Boolean Quire::op_Equality(Quire,Quire).0._State_4\, 
        \Boolean Quire::op_Equality(Quire,Quire).0._State_5\, 
        \Boolean Quire::op_Equality(Quire,Quire).0._State_6\, 
        \Boolean Quire::op_Equality(Quire,Quire).0._State_7\, 
        \Boolean Quire::op_Equality(Quire,Quire).0._State_8\);
    
    Signal \Boolean Quire::op_Equality(Quire,Quire).0._Finished\: boolean := false;
    Signal \Boolean Quire::op_Equality(Quire,Quire).0.return\: boolean := false;
    Signal \Boolean Quire::op_Equality(Quire,Quire).0.left.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Boolean Quire::op_Equality(Quire,Quire).0.right.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Boolean Quire::op_Equality(Quire,Quire).0._Started\: boolean := false;
    Signal \Boolean Quire::op_Equality(Quire,Quire).0.left.parameter.In\: \Lombiq.Arithmetics.Quire\;
    Signal \Boolean Quire::op_Equality(Quire,Quire).0.right.parameter.In\: \Lombiq.Arithmetics.Quire\;
    


    
    
    type \Quire Quire::op_RightShift(Quire,Int32).0._States\ is (
        \Quire Quire::op_RightShift(Quire,Int32).0._State_0\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_1\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_2\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_3\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_4\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_5\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_6\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_7\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_8\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_9\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_10\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_11\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_12\);
    
    Signal \Quire Quire::op_RightShift(Quire,Int32).0._Finished\: boolean := false;
    Signal \Quire Quire::op_RightShift(Quire,Int32).0.return\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_RightShift(Quire,Int32).0.left.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
    Signal \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\: boolean := false;
    Signal \Quire Quire::op_RightShift(Quire,Int32).0._Started\: boolean := false;
    Signal \Quire Quire::op_RightShift(Quire,Int32).0.left.parameter.In\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_RightShift(Quire,Int32).0.right.parameter.In\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
    Signal \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\: boolean := false;
    


    
    
    type \Quire Quire::op_LeftShift(Quire,Int32).0._States\ is (
        \Quire Quire::op_LeftShift(Quire,Int32).0._State_0\, 
        \Quire Quire::op_LeftShift(Quire,Int32).0._State_1\, 
        \Quire Quire::op_LeftShift(Quire,Int32).0._State_2\, 
        \Quire Quire::op_LeftShift(Quire,Int32).0._State_3\, 
        \Quire Quire::op_LeftShift(Quire,Int32).0._State_4\, 
        \Quire Quire::op_LeftShift(Quire,Int32).0._State_5\, 
        \Quire Quire::op_LeftShift(Quire,Int32).0._State_6\, 
        \Quire Quire::op_LeftShift(Quire,Int32).0._State_7\, 
        \Quire Quire::op_LeftShift(Quire,Int32).0._State_8\, 
        \Quire Quire::op_LeftShift(Quire,Int32).0._State_9\, 
        \Quire Quire::op_LeftShift(Quire,Int32).0._State_10\);
    
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0._Finished\: boolean := false;
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0.return\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0.left.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\: boolean := false;
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0._Started\: boolean := false;
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0.left.parameter.In\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0.right.parameter.In\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\: boolean := false;
    


    
    
    type \UInt64 Quire::op_Explicit(Quire).0._States\ is (
        \UInt64 Quire::op_Explicit(Quire).0._State_0\, 
        \UInt64 Quire::op_Explicit(Quire).0._State_1\, 
        \UInt64 Quire::op_Explicit(Quire).0._State_2\);
    
    Signal \UInt64 Quire::op_Explicit(Quire).0._Finished\: boolean := false;
    Signal \UInt64 Quire::op_Explicit(Quire).0.return\: unsigned(63 downto 0) := to_unsigned(0, 64);
    Signal \UInt64 Quire::op_Explicit(Quire).0.x.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \UInt64 Quire::op_Explicit(Quire).0._Started\: boolean := false;
    Signal \UInt64 Quire::op_Explicit(Quire).0.x.parameter.In\: \Lombiq.Arithmetics.Quire\;
    


    
    
    type \UInt32 Quire::op_Explicit(Quire).0._States\ is (
        \UInt32 Quire::op_Explicit(Quire).0._State_0\, 
        \UInt32 Quire::op_Explicit(Quire).0._State_1\, 
        \UInt32 Quire::op_Explicit(Quire).0._State_2\);
    
    Signal \UInt32 Quire::op_Explicit(Quire).0._Finished\: boolean := false;
    Signal \UInt32 Quire::op_Explicit(Quire).0.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \UInt32 Quire::op_Explicit(Quire).0.x.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \UInt32 Quire::op_Explicit(Quire).0._Started\: boolean := false;
    Signal \UInt32 Quire::op_Explicit(Quire).0.x.parameter.In\: \Lombiq.Arithmetics.Quire\;
    


    
    
    Signal \FinishedInternal\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().Posit32FusedCalculator::CalculateFusedSum(SimpleMemory)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().Posit32FusedCalculator::CalculateFusedSum(SimpleMemory)._Finished.0\: boolean := false;
    


    
    type \InternalInvocationProxy_boolean_Array\ is array (integer range <>) of boolean;
    type \Hast::InternalInvocationProxy()._RunningStates\ is (
        WaitingForStarted, 
        WaitingForFinished, 
        AfterFinished);
    

begin 

    
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._StateMachine\: process (\Clock\) 
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\: \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._States\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_0\;
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.dataIn.0\: std_logic_vector(31 downto 0) := (others => '0');
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.array\: \Lombiq.Arithmetics.Posit32_Array\(0 to 159);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.quire\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectde41e31d213f26bcb14dc4059ca0ea22b32147dbfb27f3d69d5ff482204eea98\: \Lombiq.Arithmetics.Posit32\;
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.return.0\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.3\: signed(63 downto 0) := to_signed(0, 64);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.4\: boolean := false;
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.5\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num3\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.6\: boolean := false;
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.7\: boolean := false;
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.8\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.9\: signed(63 downto 0) := to_signed(0, 64);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.10\: boolean := false;
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.11\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.12\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.13\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.dataIn.1\: std_logic_vector(31 downto 0) := (others => '0');
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.14\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.return.1\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.15\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectffd9139c321969eb0a42e1e3ae043fc0d22d96a54e32c2dc05d540c7e97af68e\: \Lombiq.Arithmetics.Posit32\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._Finished\ <= false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.DataOut\ <= (others => '0');
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).value.parameter.Out.0\ <= to_signed(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Started.0\ <= false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Started.0\ <= false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).bits.parameter.Out.0\ <= to_unsigned(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).fromBitMask.parameter.Out.0\ <= false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean)._Started.0\ <= false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire)._Started.0\ <= false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire)._Started.0\ <= false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_0\;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num\ := to_unsigned(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.dataIn.0\ := (others => '0');
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num2\ := to_unsigned(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.0\ := to_unsigned(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.1\ := to_unsigned(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.1\ := to_signed(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.2\ := to_unsigned(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.3\ := to_signed(0, 64);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.4\ := false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.5\ := to_unsigned(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num3\ := to_signed(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.6\ := false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\ := to_signed(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.7\ := false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.8\ := to_signed(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.9\ := to_signed(0, 64);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.10\ := false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.11\ := to_signed(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.12\ := to_signed(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.13\ := to_signed(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.dataIn.1\ := (others => '0');
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.14\ := to_signed(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.15\ := to_signed(0, 32);
            else 
                case \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ is 
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_0\ => 
                        
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._Started\ = true) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_2\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_1\ => 
                        
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._Started\ = true) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._Finished\ <= true;
                        else 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._Finished\ <= false;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_0\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_2\ => 
                        
                        
                        
                        
                        
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.ReadEnable\ <= true;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_3\;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_3\ => 
                        
                        if (\ReadsDone\ = true) then 
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.dataIn.0\ := \DataIn\;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num\ := ConvertStdLogicVectorToUInt32(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.dataIn.0\);
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectde41e31d213f26bcb14dc4059ca0ea22b32147dbfb27f3d69d5ff482204eea98\.\IsNull\ := false;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectde41e31d213f26bcb14dc4059ca0ea22b32147dbfb27f3d69d5ff482204eea98\.\PositBits\ := to_unsigned(0, 32);
                            
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).this.parameter.Out.0\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectde41e31d213f26bcb14dc4059ca0ea22b32147dbfb27f3d69d5ff482204eea98\;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).value.parameter.Out.0\ <= to_signed(0, 32);
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Started.0\ <= true;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_4\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_4\ => 
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Started.0\ = \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Finished.0\) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Started.0\ <= false;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectde41e31d213f26bcb14dc4059ca0ea22b32147dbfb27f3d69d5ff482204eea98\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).this.parameter.In.0\;
                            
                            
                            
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32).x.parameter.Out.0\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectde41e31d213f26bcb14dc4059ca0ea22b32147dbfb27f3d69d5ff482204eea98\;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Started.0\ <= true;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_5\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_5\ => 
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Started.0\ = \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Started.0\ <= false;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.return.0\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32).return.0\;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.quire\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.return.0\;
                            
                            
                            
                            
                            
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_6\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_6\ => 
                        
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(8, 32)) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_7\;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.0\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.0\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num\ / to_unsigned(160, 32);
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_7\ => 
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num2\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.0\;
                        
                        
                        
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_8\;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_8\ => 
                        
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.1\ >= to_signed(8, 32)) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_9\;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.1\ := to_signed(0, 32);
                        else 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.1\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.1\ + to_signed(1, 32);
                        end if;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.1\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num\ / to_unsigned(160, 32);
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_9\ => 
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.2\ := SmartResize(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.1\ * to_unsigned(160, 32), 32);
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.3\ := signed(SmartResize(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num\ - \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.2\, 64));
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_10\;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_10\ => 
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.4\ := (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.3\) /= to_signed(0, 64);

                        
                        
                        

                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.4\) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_12\;
                        else 
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_11\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_11\ => 
                        
                        
                        
                        
                        
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num3\ := to_signed(0, 32);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_13\;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_12\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.5\ := SmartResize(unsigned(signed(SmartResize((\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num2\), 64)) + to_signed(1, 64)), 32);
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num2\ := (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.5\);
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ = \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_12\) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_11\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_13\ => 
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.6\ := SmartResize((\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num3\), 64) < signed(SmartResize((\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num2\), 64));
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.6\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\ := to_signed(0, 32);
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_15\;
                        else 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_14\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_14\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectffd9139c321969eb0a42e1e3ae043fc0d22d96a54e32c2dc05d540c7e97af68e\.\IsNull\ := false;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectffd9139c321969eb0a42e1e3ae043fc0d22d96a54e32c2dc05d540c7e97af68e\.\PositBits\ := to_unsigned(0, 32);
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).this.parameter.Out.0\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectffd9139c321969eb0a42e1e3ae043fc0d22d96a54e32c2dc05d540c7e97af68e\;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).q.parameter.Out.0\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.quire\;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire)._Started.0\ <= true;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_27\;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_15\ => 
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.7\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\ < to_signed(160, 32);
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.7\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.8\ := SmartResize(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num3\ * to_signed(160, 32), 32);
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_17\;
                        else 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_16\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_16\ => 
                        
                        
                        
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).posits.parameter.Out.0\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.array\;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).startingValue.parameter.Out.0\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.quire\;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire)._Started.0\ <= true;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_26\;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_17\ => 
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.9\ := SmartResize(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.8\ + \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\, 64);
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_18\;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_18\ => 
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.10\ := (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.9\) < signed(SmartResize((\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num\), 64));

                        
                        
                        
                        

                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.10\) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_20\;
                        else 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_24\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_19\ => 
                        
                        
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.14\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\ + to_signed(1, 32);
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.14\;
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ = \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_19\) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_15\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_20\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.array\(to_integer(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\)).\IsNull\ := false;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.array\(to_integer(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\)).\PositBits\ := to_unsigned(0, 32);
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.11\ := SmartResize(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num3\ * to_signed(160, 32), 32);
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.12\ := to_signed(1, 32) + \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.11\;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_21\;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_21\ => 
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.13\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.12\ + \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\;
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.CellIndex\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.13\;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.ReadEnable\ <= true;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_22\;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_22\ => 
                        
                        if (\ReadsDone\ = true) then 
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.dataIn.1\ := \DataIn\;
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).this.parameter.Out.0\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.array\(to_integer(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\));
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).bits.parameter.Out.0\ <= ConvertStdLogicVectorToUInt32(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.dataIn.1\);
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).fromBitMask.parameter.Out.0\ <= true;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean)._Started.0\ <= true;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_23\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_23\ => 
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean)._Started.0\ = \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean)._Finished.0\) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean)._Started.0\ <= false;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.array\(to_integer(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\)) := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).this.parameter.In.0\;
                            
                            if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ = \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_23\) then 
                                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_19\;
                            end if;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_24\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.array\(to_integer(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\)).\IsNull\ := false;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.array\(to_integer(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\)).\PositBits\ := to_unsigned(0, 32);
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).this.parameter.Out.0\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.array\(to_integer(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\));
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).value.parameter.Out.0\ <= to_signed(0, 32);
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Started.0\ <= true;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_25\;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_25\ => 
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Started.0\ = \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Finished.0\) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Started.0\ <= false;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.array\(to_integer(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\)) := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).this.parameter.In.0\;
                            
                            if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ = \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_25\) then 
                                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_19\;
                            end if;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_26\ => 
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire)._Started.0\ = \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire)._Finished.0\) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire)._Started.0\ <= false;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.return.1\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).return.0\;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.array\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).posits.parameter.In.0\;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.quire\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).startingValue.parameter.In.0\;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.quire\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.return.1\;
                            
                            
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.15\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num3\ + to_signed(1, 32);
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num3\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.15\;
                            
                            if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ = \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_26\) then 
                                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_13\;
                            end if;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_27\ => 
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire)._Started.0\ = \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire)._Finished.0\) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire)._Started.0\ <= false;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectffd9139c321969eb0a42e1e3ae043fc0d22d96a54e32c2dc05d540c7e97af68e\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).this.parameter.In.0\;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.quire\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).q.parameter.In.0\;
                            
                            
                            
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.WriteEnable\ <= true;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.DataOut\ <= ConvertUInt32ToStdLogicVector(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectffd9139c321969eb0a42e1e3ae043fc0d22d96a54e32c2dc05d540c7e97af68e\.\PositBits\);
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_28\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_28\ => 
                        
                        if (\WritesDone\ = true) then 
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_1\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::.ctor(UInt32,Boolean).0._StateMachine\: process (\Clock\) 
        Variable \Posit32::.ctor(UInt32,Boolean).0._State\: \Posit32::.ctor(UInt32,Boolean).0._States\ := \Posit32::.ctor(UInt32,Boolean).0._State_0\;
        Variable \Posit32::.ctor(UInt32,Boolean).0.this\: \Lombiq.Arithmetics.Posit32\;
        Variable \Posit32::.ctor(UInt32,Boolean).0.bits\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::.ctor(UInt32,Boolean).0.fromBitMask\: boolean := false;
        Variable \Posit32::.ctor(UInt32,Boolean).0.conditional07306ef17ce6eacdbdd521687c7db8bbabd2dc9ca02b65fce7cdbd581ebb7be6\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::.ctor(UInt32,Boolean).0._Finished\ <= false;
                \Posit32::.ctor(UInt32,Boolean).0._State\ := \Posit32::.ctor(UInt32,Boolean).0._State_0\;
                \Posit32::.ctor(UInt32,Boolean).0.bits\ := to_unsigned(0, 32);
                \Posit32::.ctor(UInt32,Boolean).0.fromBitMask\ := false;
                \Posit32::.ctor(UInt32,Boolean).0.conditional07306ef17ce6eacdbdd521687c7db8bbabd2dc9ca02b65fce7cdbd581ebb7be6\ := to_unsigned(0, 32);
            else 
                case \Posit32::.ctor(UInt32,Boolean).0._State\ is 
                    when \Posit32::.ctor(UInt32,Boolean).0._State_0\ => 
                        
                        
                        if (\Posit32::.ctor(UInt32,Boolean).0._Started\ = true) then 
                            \Posit32::.ctor(UInt32,Boolean).0._State\ := \Posit32::.ctor(UInt32,Boolean).0._State_2\;
                        end if;
                        
                    when \Posit32::.ctor(UInt32,Boolean).0._State_1\ => 
                        
                        
                        if (\Posit32::.ctor(UInt32,Boolean).0._Started\ = true) then 
                            \Posit32::.ctor(UInt32,Boolean).0._Finished\ <= true;
                        else 
                            \Posit32::.ctor(UInt32,Boolean).0._Finished\ <= false;
                            \Posit32::.ctor(UInt32,Boolean).0._State\ := \Posit32::.ctor(UInt32,Boolean).0._State_0\;
                        end if;
                        
                        \Posit32::.ctor(UInt32,Boolean).0.this.parameter.Out\ <= \Posit32::.ctor(UInt32,Boolean).0.this\;
                        
                    when \Posit32::.ctor(UInt32,Boolean).0._State_2\ => 
                        \Posit32::.ctor(UInt32,Boolean).0.this\ := \Posit32::.ctor(UInt32,Boolean).0.this.parameter.In\;
                        \Posit32::.ctor(UInt32,Boolean).0.bits\ := \Posit32::.ctor(UInt32,Boolean).0.bits.parameter.In\;
                        \Posit32::.ctor(UInt32,Boolean).0.fromBitMask\ := \Posit32::.ctor(UInt32,Boolean).0.fromBitMask.parameter.In\;
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(UInt32,Boolean).0.conditional07306ef17ce6eacdbdd521687c7db8bbabd2dc9ca02b65fce7cdbd581ebb7be6\ := \Posit32::.ctor(UInt32,Boolean).0.bits\;
                        
                        
                        
                        \Posit32::.ctor(UInt32,Boolean).0.this\.\PositBits\ := (\Posit32::.ctor(UInt32,Boolean).0.conditional07306ef17ce6eacdbdd521687c7db8bbabd2dc9ca02b65fce7cdbd581ebb7be6\);
                        \Posit32::.ctor(UInt32,Boolean).0._State\ := \Posit32::.ctor(UInt32,Boolean).0._State_1\;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::.ctor(Quire).0._StateMachine\: process (\Clock\) 
        Variable \Posit32::.ctor(Quire).0._State\: \Posit32::.ctor(Quire).0._States\ := \Posit32::.ctor(Quire).0._State_0\;
        Variable \Posit32::.ctor(Quire).0.this\: \Lombiq.Arithmetics.Posit32\;
        Variable \Posit32::.ctor(Quire).0.q\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::.ctor(Quire).0.signBit\: boolean := false;
        Variable \Posit32::.ctor(Quire).0.num\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::.ctor(Quire).0.num2\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Posit32::.ctor(Quire).0.return.0\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::.ctor(Quire).0.return.1\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.0\: boolean := false;
        Variable \Posit32::.ctor(Quire).0.return.2\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::.ctor(Quire).0.return.3\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::.ctor(Quire).0.return.4\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::.ctor(Quire).0.return.5\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.1\: boolean := false;
        Variable \Posit32::.ctor(Quire).0.return.6\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::.ctor(Quire).0.return.7\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::.ctor(Quire).0.return.8\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Posit32::.ctor(Quire).0.num3\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.3\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.4\: boolean := false;
        Variable \Posit32::.ctor(Quire).0.num4\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.5\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::.ctor(Quire).0.num5\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.6\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.7\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.8\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.9\: boolean := false;
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.10\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.11\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::.ctor(Quire).0.return.9\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::.ctor(Quire).0.return.10\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::.ctor(Quire).0.return.11\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::.ctor(Quire).0._Finished\ <= false;
                \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).right.parameter.Out.0\ <= to_signed(0, 32);
                \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ <= false;
                \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\ <= false;
                \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire)._Started.0\ <= false;
                \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).right.parameter.Out.0\ <= to_unsigned(0, 32);
                \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32)._Started.0\ <= false;
                \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\ <= to_signed(0, 32);
                \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ <= false;
                \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire)._Started.0\ <= false;
                \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).signBit.parameter.Out.0\ <= false;
                \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).regimeKValue.parameter.Out.0\ <= to_signed(0, 32);
                \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).exponentBits.parameter.Out.0\ <= to_unsigned(0, 32);
                \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).fractionBits.parameter.Out.0\ <= to_unsigned(0, 32);
                \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32)._Started.0\ <= false;
                \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_0\;
                \Posit32::.ctor(Quire).0.signBit\ := false;
                \Posit32::.ctor(Quire).0.num\ := to_signed(0, 32);
                \Posit32::.ctor(Quire).0.num2\ := to_unsigned(0, 64);
                \Posit32::.ctor(Quire).0.return.1\ := to_unsigned(0, 64);
                \Posit32::.ctor(Quire).0.binaryOperationResult.0\ := false;
                \Posit32::.ctor(Quire).0.return.5\ := to_unsigned(0, 64);
                \Posit32::.ctor(Quire).0.binaryOperationResult.1\ := false;
                \Posit32::.ctor(Quire).0.binaryOperationResult.2\ := to_signed(0, 32);
                \Posit32::.ctor(Quire).0.return.8\ := to_unsigned(0, 64);
                \Posit32::.ctor(Quire).0.num3\ := to_signed(0, 32);
                \Posit32::.ctor(Quire).0.binaryOperationResult.3\ := to_signed(0, 32);
                \Posit32::.ctor(Quire).0.binaryOperationResult.4\ := false;
                \Posit32::.ctor(Quire).0.num4\ := to_signed(0, 32);
                \Posit32::.ctor(Quire).0.binaryOperationResult.5\ := to_signed(0, 32);
                \Posit32::.ctor(Quire).0.num5\ := to_unsigned(0, 32);
                \Posit32::.ctor(Quire).0.binaryOperationResult.6\ := to_signed(0, 32);
                \Posit32::.ctor(Quire).0.binaryOperationResult.7\ := to_signed(0, 32);
                \Posit32::.ctor(Quire).0.binaryOperationResult.8\ := to_unsigned(0, 32);
                \Posit32::.ctor(Quire).0.binaryOperationResult.9\ := false;
                \Posit32::.ctor(Quire).0.binaryOperationResult.10\ := to_signed(0, 32);
                \Posit32::.ctor(Quire).0.binaryOperationResult.11\ := to_unsigned(0, 32);
                \Posit32::.ctor(Quire).0.return.10\ := to_unsigned(0, 32);
                \Posit32::.ctor(Quire).0.return.11\ := to_unsigned(0, 32);
            else 
                case \Posit32::.ctor(Quire).0._State\ is 
                    when \Posit32::.ctor(Quire).0._State_0\ => 
                        
                        
                        if (\Posit32::.ctor(Quire).0._Started\ = true) then 
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_2\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_1\ => 
                        
                        
                        if (\Posit32::.ctor(Quire).0._Started\ = true) then 
                            \Posit32::.ctor(Quire).0._Finished\ <= true;
                        else 
                            \Posit32::.ctor(Quire).0._Finished\ <= false;
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_0\;
                        end if;
                        
                        \Posit32::.ctor(Quire).0.this.parameter.Out\ <= \Posit32::.ctor(Quire).0.this\;
                        \Posit32::.ctor(Quire).0.q.parameter.Out\ <= \Posit32::.ctor(Quire).0.q\;
                        
                    when \Posit32::.ctor(Quire).0._State_2\ => 
                        \Posit32::.ctor(Quire).0.this\ := \Posit32::.ctor(Quire).0.this.parameter.In\;
                        \Posit32::.ctor(Quire).0.q\ := \Posit32::.ctor(Quire).0.q.parameter.In\;
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.this\.\PositBits\ := "10000000000000000000000000000000";
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.signBit\ := false;
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.num\ := to_signed(511, 32);
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.q\;
                        \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).right.parameter.Out.0\ <= to_signed(448, 32);
                        \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ <= true;
                        \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_3\;
                        
                    when \Posit32::.ctor(Quire).0._State_3\ => 
                        
                        if (\Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ = \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.0\ := \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).return.0\;
                            \Posit32::.ctor(Quire).0.q\ := \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.In.0\;
                            
                            \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).x.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.return.0\;
                            \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\ <= true;
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_4\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_4\ => 
                        
                        if (\Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\ = \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.1\ := \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).return.0\;
                            \Posit32::.ctor(Quire).0.return.0\ := \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).x.parameter.In.0\;
                            \Posit32::.ctor(Quire).0.num2\ := \Posit32::.ctor(Quire).0.return.1\;
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32::.ctor(Quire).0.binaryOperationResult.0\ := \Posit32::.ctor(Quire).0.num2\ >= "1000000000000000000000000000000000000000000000000000000000000000";

                            
                            
                            

                            if (\Posit32::.ctor(Quire).0.binaryOperationResult.0\) then 
                                \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_6\;
                            else 
                                
                                \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_5\;
                            end if;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_5\ => 
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.q\;
                        \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).right.parameter.Out.0\ <= to_signed(448, 32);
                        \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ <= true;
                        \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_9\;
                        
                    when \Posit32::.ctor(Quire).0._State_6\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire).q.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.q\;
                        \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire)._Started.0\ <= true;
                        \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_7\;
                        
                    when \Posit32::.ctor(Quire).0._State_7\ => 
                        
                        if (\Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire)._Started.0\ = \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.2\ := \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire).return.0\;
                            \Posit32::.ctor(Quire).0.q\ := \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire).q.parameter.In.0\;
                            \Posit32::.ctor(Quire).0.q\ := \Posit32::.ctor(Quire).0.return.2\;
                            
                            
                            
                            
                            \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).left.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.q\;
                            \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).right.parameter.Out.0\ <= to_unsigned(1, 32);
                            \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32)._Started.0\ <= true;
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_8\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_8\ => 
                        
                        if (\Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32)._Started.0\ = \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.3\ := \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).return.0\;
                            \Posit32::.ctor(Quire).0.q\ := \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).left.parameter.In.0\;
                            \Posit32::.ctor(Quire).0.q\ := \Posit32::.ctor(Quire).0.return.3\;
                            
                            
                            
                            \Posit32::.ctor(Quire).0.signBit\ := true;
                            
                            if (\Posit32::.ctor(Quire).0._State\ = \Posit32::.ctor(Quire).0._State_8\) then 
                                \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_5\;
                            end if;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_9\ => 
                        
                        if (\Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ = \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.4\ := \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).return.0\;
                            \Posit32::.ctor(Quire).0.q\ := \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.In.0\;
                            
                            \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).x.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.return.4\;
                            \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\ <= true;
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_10\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_10\ => 
                        
                        if (\Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\ = \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.5\ := \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).return.0\;
                            \Posit32::.ctor(Quire).0.return.4\ := \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).x.parameter.In.0\;
                            \Posit32::.ctor(Quire).0.num2\ := \Posit32::.ctor(Quire).0.return.5\;
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_11\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_11\ => 
                        
                        
                        
                        \Posit32::.ctor(Quire).0.binaryOperationResult.1\ := \Posit32::.ctor(Quire).0.num2\ < "1000000000000000000000000000000000000000000000000000000000000000";
                        if (\Posit32::.ctor(Quire).0.binaryOperationResult.1\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.q\;
                            \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\ <= to_signed(1, 32);
                            \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ <= true;
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_13\;
                        else 
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_12\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_12\ => 
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.binaryOperationResult.3\ := \Posit32::.ctor(Quire).0.num\ - to_signed(240, 32);
                        \Posit32::.ctor(Quire).0.num3\ := \Posit32::.ctor(Quire).0.binaryOperationResult.3\;
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.binaryOperationResult.4\ := \Posit32::.ctor(Quire).0.num\ = to_signed(0, 32);

                        
                        
                        

                        if (\Posit32::.ctor(Quire).0.binaryOperationResult.4\) then 
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_17\;
                        else 
                            
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_16\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_13\ => 
                        
                        if (\Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ = \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.6\ := \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).return.0\;
                            \Posit32::.ctor(Quire).0.q\ := \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.In.0\;
                            \Posit32::.ctor(Quire).0.q\ := \Posit32::.ctor(Quire).0.return.6\;
                            
                            
                            
                            \Posit32::.ctor(Quire).0.binaryOperationResult.2\ := \Posit32::.ctor(Quire).0.num\ - to_signed(1, 32);
                            \Posit32::.ctor(Quire).0.num\ := \Posit32::.ctor(Quire).0.binaryOperationResult.2\;
                            
                            
                            
                            
                            \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.q\;
                            \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).right.parameter.Out.0\ <= to_signed(448, 32);
                            \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ <= true;
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_14\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_14\ => 
                        
                        if (\Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ = \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.7\ := \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).return.0\;
                            \Posit32::.ctor(Quire).0.q\ := \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.In.0\;
                            
                            \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).x.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.return.7\;
                            \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\ <= true;
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_15\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_15\ => 
                        
                        if (\Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\ = \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.8\ := \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).return.0\;
                            \Posit32::.ctor(Quire).0.return.7\ := \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).x.parameter.In.0\;
                            \Posit32::.ctor(Quire).0.num2\ := \Posit32::.ctor(Quire).0.return.8\;
                            
                            if (\Posit32::.ctor(Quire).0._State\ = \Posit32::.ctor(Quire).0._State_15\) then 
                                \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_11\;
                            end if;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_16\ => 
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.binaryOperationResult.5\ := \Posit32::.ctor(Quire).0.num3\ / to_signed(4, 32);
                        \Posit32::.ctor(Quire).0.num4\ := \Posit32::.ctor(Quire).0.binaryOperationResult.5\;
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.binaryOperationResult.6\ := \Posit32::.ctor(Quire).0.num3\ / to_signed(4, 32);
                        \Posit32::.ctor(Quire).0.binaryOperationResult.7\ := SmartResize(\Posit32::.ctor(Quire).0.binaryOperationResult.6\ * to_signed(4, 32), 32);
                        \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_18\;
                        
                    when \Posit32::.ctor(Quire).0._State_17\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.this\.\PositBits\ := to_unsigned(0, 32);
                        
                        
                        
                        \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_1\;
                        
                        if (\Posit32::.ctor(Quire).0._State\ = \Posit32::.ctor(Quire).0._State_17\) then 
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_16\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_18\ => 
                        
                        \Posit32::.ctor(Quire).0.binaryOperationResult.8\ := unsigned(\Posit32::.ctor(Quire).0.num3\ - \Posit32::.ctor(Quire).0.binaryOperationResult.7\);
                        \Posit32::.ctor(Quire).0.num5\ := (\Posit32::.ctor(Quire).0.binaryOperationResult.8\);
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_19\;
                        
                    when \Posit32::.ctor(Quire).0._State_19\ => 
                        
                        \Posit32::.ctor(Quire).0.binaryOperationResult.9\ := signed(SmartResize((\Posit32::.ctor(Quire).0.num5\), 64)) < to_signed(0, 64);

                        
                        
                        

                        if (\Posit32::.ctor(Quire).0.binaryOperationResult.9\) then 
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_21\;
                        else 
                            
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_20\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_20\ => 
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.q\;
                        \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).right.parameter.Out.0\ <= to_signed(480, 32);
                        \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ <= true;
                        \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_22\;
                        
                    when \Posit32::.ctor(Quire).0._State_21\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.binaryOperationResult.10\ := \Posit32::.ctor(Quire).0.num4\ - to_signed(1, 32);
                        \Posit32::.ctor(Quire).0.num4\ := \Posit32::.ctor(Quire).0.binaryOperationResult.10\;
                        
                        
                        
                        \Posit32::.ctor(Quire).0.binaryOperationResult.11\ := SmartResize(unsigned(signed(SmartResize((\Posit32::.ctor(Quire).0.num5\), 64)) + to_signed(4, 64)), 32);
                        \Posit32::.ctor(Quire).0.num5\ := (\Posit32::.ctor(Quire).0.binaryOperationResult.11\);
                        
                        if (\Posit32::.ctor(Quire).0._State\ = \Posit32::.ctor(Quire).0._State_21\) then 
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_20\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_22\ => 
                        
                        if (\Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ = \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.9\ := \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).return.0\;
                            \Posit32::.ctor(Quire).0.q\ := \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.In.0\;
                            
                            \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire).x.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.return.9\;
                            \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire)._Started.0\ <= true;
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_23\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_23\ => 
                        
                        if (\Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire)._Started.0\ = \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.10\ := \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire).return.0\;
                            \Posit32::.ctor(Quire).0.return.9\ := \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire).x.parameter.In.0\;
                            
                            \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).signBit.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.signBit\;
                            \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).regimeKValue.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.num4\;
                            \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).exponentBits.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.num5\;
                            \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).fractionBits.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.return.10\;
                            \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32)._Started.0\ <= true;
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_24\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_24\ => 
                        
                        if (\Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32)._Started.0\ = \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.11\ := \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).return.0\;
                            \Posit32::.ctor(Quire).0.this\.\PositBits\ := \Posit32::.ctor(Quire).0.return.11\;
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_1\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::.ctor(UInt32).0._StateMachine\: process (\Clock\) 
        Variable \Posit32::.ctor(UInt32).0._State\: \Posit32::.ctor(UInt32).0._States\ := \Posit32::.ctor(UInt32).0._State_0\;
        Variable \Posit32::.ctor(UInt32).0.this\: \Lombiq.Arithmetics.Posit32\;
        Variable \Posit32::.ctor(UInt32).0.value\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::.ctor(UInt32).0._Finished\ <= false;
                \Posit32::.ctor(UInt32).0._State\ := \Posit32::.ctor(UInt32).0._State_0\;
                \Posit32::.ctor(UInt32).0.value\ := to_unsigned(0, 32);
            else 
                case \Posit32::.ctor(UInt32).0._State\ is 
                    when \Posit32::.ctor(UInt32).0._State_0\ => 
                        
                        
                        if (\Posit32::.ctor(UInt32).0._Started\ = true) then 
                            \Posit32::.ctor(UInt32).0._State\ := \Posit32::.ctor(UInt32).0._State_2\;
                        end if;
                        
                    when \Posit32::.ctor(UInt32).0._State_1\ => 
                        
                        
                        if (\Posit32::.ctor(UInt32).0._Started\ = true) then 
                            \Posit32::.ctor(UInt32).0._Finished\ <= true;
                        else 
                            \Posit32::.ctor(UInt32).0._Finished\ <= false;
                            \Posit32::.ctor(UInt32).0._State\ := \Posit32::.ctor(UInt32).0._State_0\;
                        end if;
                        
                        \Posit32::.ctor(UInt32).0.this.parameter.Out\ <= \Posit32::.ctor(UInt32).0.this\;
                        
                    when \Posit32::.ctor(UInt32).0._State_2\ => 
                        \Posit32::.ctor(UInt32).0.this\ := \Posit32::.ctor(UInt32).0.this.parameter.In\;
                        \Posit32::.ctor(UInt32).0.value\ := \Posit32::.ctor(UInt32).0.value.parameter.In\;
                        
                        
                        
                        \Posit32::.ctor(UInt32).0.this\.\PositBits\ := to_unsigned(0, 32);
                        \Posit32::.ctor(UInt32).0._State\ := \Posit32::.ctor(UInt32).0._State_1\;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::.ctor(Int32).0._StateMachine\: process (\Clock\) 
        Variable \Posit32::.ctor(Int32).0._State\: \Posit32::.ctor(Int32).0._States\ := \Posit32::.ctor(Int32).0._State_0\;
        Variable \Posit32::.ctor(Int32).0.this\: \Lombiq.Arithmetics.Posit32\;
        Variable \Posit32::.ctor(Int32).0.value\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::.ctor(Int32).0.conditional2430432b7cbc58715e662a8c82abb8a42239e5b92d4c7ea6c2c87a87483f3331\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::.ctor(Int32).0.object62f645adbfb4d116e9dadbde41fc03ee8eecadf80abd12f7fbc8d9dfa7162321\: \Lombiq.Arithmetics.Posit32\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::.ctor(Int32).0._Finished\ <= false;
                \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32).value.parameter.Out.0\ <= to_unsigned(0, 32);
                \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32)._Started.0\ <= false;
                \Posit32::.ctor(Int32).0._State\ := \Posit32::.ctor(Int32).0._State_0\;
                \Posit32::.ctor(Int32).0.value\ := to_signed(0, 32);
                \Posit32::.ctor(Int32).0.conditional2430432b7cbc58715e662a8c82abb8a42239e5b92d4c7ea6c2c87a87483f3331\ := to_unsigned(0, 32);
            else 
                case \Posit32::.ctor(Int32).0._State\ is 
                    when \Posit32::.ctor(Int32).0._State_0\ => 
                        
                        
                        if (\Posit32::.ctor(Int32).0._Started\ = true) then 
                            \Posit32::.ctor(Int32).0._State\ := \Posit32::.ctor(Int32).0._State_2\;
                        end if;
                        
                    when \Posit32::.ctor(Int32).0._State_1\ => 
                        
                        
                        if (\Posit32::.ctor(Int32).0._Started\ = true) then 
                            \Posit32::.ctor(Int32).0._Finished\ <= true;
                        else 
                            \Posit32::.ctor(Int32).0._Finished\ <= false;
                            \Posit32::.ctor(Int32).0._State\ := \Posit32::.ctor(Int32).0._State_0\;
                        end if;
                        
                        \Posit32::.ctor(Int32).0.this.parameter.Out\ <= \Posit32::.ctor(Int32).0.this\;
                        
                    when \Posit32::.ctor(Int32).0._State_2\ => 
                        \Posit32::.ctor(Int32).0.this\ := \Posit32::.ctor(Int32).0.this.parameter.In\;
                        \Posit32::.ctor(Int32).0.value\ := \Posit32::.ctor(Int32).0.value.parameter.In\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Int32).0.object62f645adbfb4d116e9dadbde41fc03ee8eecadf80abd12f7fbc8d9dfa7162321\.\IsNull\ := false;
                        \Posit32::.ctor(Int32).0.object62f645adbfb4d116e9dadbde41fc03ee8eecadf80abd12f7fbc8d9dfa7162321\.\PositBits\ := to_unsigned(0, 32);
                        
                        
                        \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32).this.parameter.Out.0\ <= \Posit32::.ctor(Int32).0.object62f645adbfb4d116e9dadbde41fc03ee8eecadf80abd12f7fbc8d9dfa7162321\;
                        \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32).value.parameter.Out.0\ <= to_unsigned(0, 32);
                        \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32)._Started.0\ <= true;
                        \Posit32::.ctor(Int32).0._State\ := \Posit32::.ctor(Int32).0._State_3\;
                        
                    when \Posit32::.ctor(Int32).0._State_3\ => 
                        
                        if (\Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32)._Started.0\ = \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32)._Finished.0\) then 
                            \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32)._Started.0\ <= false;
                            \Posit32::.ctor(Int32).0.object62f645adbfb4d116e9dadbde41fc03ee8eecadf80abd12f7fbc8d9dfa7162321\ := \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32).this.parameter.In.0\;
                            
                            
                            
                            \Posit32::.ctor(Int32).0.conditional2430432b7cbc58715e662a8c82abb8a42239e5b92d4c7ea6c2c87a87483f3331\ := to_unsigned(0, 32);
                            
                            
                            
                            \Posit32::.ctor(Int32).0.this\.\PositBits\ := to_unsigned(0, 32);
                            \Posit32::.ctor(Int32).0._State\ := \Posit32::.ctor(Int32).0._State_1\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::IsNaN().0._StateMachine\: process (\Clock\) 
        Variable \Posit32::IsNaN().0._State\: \Posit32::IsNaN().0._States\ := \Posit32::IsNaN().0._State_0\;
        Variable \Posit32::IsNaN().0.this\: \Lombiq.Arithmetics.Posit32\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::IsNaN().0._Finished\ <= false;
                \Posit32::IsNaN().0.return\ <= false;
                \Posit32::IsNaN().0._State\ := \Posit32::IsNaN().0._State_0\;
            else 
                case \Posit32::IsNaN().0._State\ is 
                    when \Posit32::IsNaN().0._State_0\ => 
                        
                        
                        if (\Posit32::IsNaN().0._Started\ = true) then 
                            \Posit32::IsNaN().0._State\ := \Posit32::IsNaN().0._State_2\;
                        end if;
                        
                    when \Posit32::IsNaN().0._State_1\ => 
                        
                        
                        if (\Posit32::IsNaN().0._Started\ = true) then 
                            \Posit32::IsNaN().0._Finished\ <= true;
                        else 
                            \Posit32::IsNaN().0._Finished\ <= false;
                            \Posit32::IsNaN().0._State\ := \Posit32::IsNaN().0._State_0\;
                        end if;
                        
                    when \Posit32::IsNaN().0._State_2\ => 
                        \Posit32::IsNaN().0.this\ := \Posit32::IsNaN().0.this.parameter.In\;
                        
                        
                        
                        \Posit32::IsNaN().0.return\ <= false;
                        \Posit32::IsNaN().0._State\ := \Posit32::IsNaN().0._State_1\;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::EncodeRegimeBits(Int32).0._StateMachine\: process (\Clock\) 
        Variable \Posit32::EncodeRegimeBits(Int32).0._State\: \Posit32::EncodeRegimeBits(Int32).0._States\ := \Posit32::EncodeRegimeBits(Int32).0._State_0\;
        Variable \Posit32::EncodeRegimeBits(Int32).0.regimeKValue\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.0\: boolean := false;
        Variable \Posit32::EncodeRegimeBits(Int32).0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::EncodeRegimeBits(Int32).0.return.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.4\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.5\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.6\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::EncodeRegimeBits(Int32).0.unaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.7\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::EncodeRegimeBits(Int32).0._Finished\ <= false;
                \Posit32::EncodeRegimeBits(Int32).0.return\ <= to_unsigned(0, 32);
                \Posit32::EncodeRegimeBits(Int32).0.Posit32::GetMostSignificantOnePosition(UInt32).bits.parameter.Out.0\ <= to_unsigned(0, 32);
                \Posit32::EncodeRegimeBits(Int32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Started.0\ <= false;
                \Posit32::EncodeRegimeBits(Int32).0._State\ := \Posit32::EncodeRegimeBits(Int32).0._State_0\;
                \Posit32::EncodeRegimeBits(Int32).0.regimeKValue\ := to_signed(0, 32);
                \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.0\ := false;
                \Posit32::EncodeRegimeBits(Int32).0.num\ := to_unsigned(0, 32);
                \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.1\ := to_signed(0, 32);
                \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.2\ := to_signed(0, 32);
                \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.3\ := to_unsigned(0, 32);
                \Posit32::EncodeRegimeBits(Int32).0.return.0\ := to_unsigned(0, 8);
                \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.4\ := to_signed(0, 32);
                \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.5\ := to_signed(0, 32);
                \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.6\ := to_unsigned(0, 32);
                \Posit32::EncodeRegimeBits(Int32).0.unaryOperationResult.0\ := to_signed(0, 32);
                \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.7\ := to_unsigned(0, 32);
            else 
                case \Posit32::EncodeRegimeBits(Int32).0._State\ is 
                    when \Posit32::EncodeRegimeBits(Int32).0._State_0\ => 
                        
                        
                        if (\Posit32::EncodeRegimeBits(Int32).0._Started\ = true) then 
                            \Posit32::EncodeRegimeBits(Int32).0._State\ := \Posit32::EncodeRegimeBits(Int32).0._State_2\;
                        end if;
                        
                    when \Posit32::EncodeRegimeBits(Int32).0._State_1\ => 
                        
                        
                        if (\Posit32::EncodeRegimeBits(Int32).0._Started\ = true) then 
                            \Posit32::EncodeRegimeBits(Int32).0._Finished\ <= true;
                        else 
                            \Posit32::EncodeRegimeBits(Int32).0._Finished\ <= false;
                            \Posit32::EncodeRegimeBits(Int32).0._State\ := \Posit32::EncodeRegimeBits(Int32).0._State_0\;
                        end if;
                        
                    when \Posit32::EncodeRegimeBits(Int32).0._State_2\ => 
                        \Posit32::EncodeRegimeBits(Int32).0.regimeKValue\ := \Posit32::EncodeRegimeBits(Int32).0.regimeKValue.parameter.In\;
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.0\ := \Posit32::EncodeRegimeBits(Int32).0.regimeKValue\ > to_signed(0, 32);

                        
                        
                        

                        if (\Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.0\) then 
                            \Posit32::EncodeRegimeBits(Int32).0._State\ := \Posit32::EncodeRegimeBits(Int32).0._State_4\;
                        else 
                            
                            \Posit32::EncodeRegimeBits(Int32).0._State\ := \Posit32::EncodeRegimeBits(Int32).0._State_3\;
                        end if;
                        
                    when \Posit32::EncodeRegimeBits(Int32).0._State_3\ => 
                        
                        
                        
                        
                        \Posit32::EncodeRegimeBits(Int32).0.unaryOperationResult.0\ := -\Posit32::EncodeRegimeBits(Int32).0.regimeKValue\;
                        \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.7\ := shift_right(to_unsigned(1073741824, 32), to_integer(unsigned(SmartResize(\Posit32::EncodeRegimeBits(Int32).0.unaryOperationResult.0\, 5) and "11111")));
                        \Posit32::EncodeRegimeBits(Int32).0.return\ <= \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.7\;
                        \Posit32::EncodeRegimeBits(Int32).0._State\ := \Posit32::EncodeRegimeBits(Int32).0._State_1\;
                        
                    when \Posit32::EncodeRegimeBits(Int32).0._State_4\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.1\ := \Posit32::EncodeRegimeBits(Int32).0.regimeKValue\ + to_signed(1, 32);
                        \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.2\ := shift_left(to_signed(1, 32), to_integer(unsigned(SmartResize(\Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.1\, 5))));
                        \Posit32::EncodeRegimeBits(Int32).0._State\ := \Posit32::EncodeRegimeBits(Int32).0._State_5\;
                        
                    when \Posit32::EncodeRegimeBits(Int32).0._State_5\ => 
                        
                        \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.3\ := unsigned((\Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.2\) - to_signed(1, 32));
                        \Posit32::EncodeRegimeBits(Int32).0.num\ := (\Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.3\);
                        
                        
                        
                        
                        \Posit32::EncodeRegimeBits(Int32).0.Posit32::GetMostSignificantOnePosition(UInt32).bits.parameter.Out.0\ <= \Posit32::EncodeRegimeBits(Int32).0.num\;
                        \Posit32::EncodeRegimeBits(Int32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Started.0\ <= true;
                        \Posit32::EncodeRegimeBits(Int32).0._State\ := \Posit32::EncodeRegimeBits(Int32).0._State_6\;
                        
                    when \Posit32::EncodeRegimeBits(Int32).0._State_6\ => 
                        
                        if (\Posit32::EncodeRegimeBits(Int32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Started.0\ = \Posit32::EncodeRegimeBits(Int32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Finished.0\) then 
                            \Posit32::EncodeRegimeBits(Int32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Started.0\ <= false;
                            \Posit32::EncodeRegimeBits(Int32).0.return.0\ := \Posit32::EncodeRegimeBits(Int32).0.Posit32::GetMostSignificantOnePosition(UInt32).return.0\;
                            \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.4\ := to_signed(32, 32) - signed(SmartResize((\Posit32::EncodeRegimeBits(Int32).0.return.0\), 32));
                            \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.5\ := \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.4\ - to_signed(1, 32);
                            \Posit32::EncodeRegimeBits(Int32).0._State\ := \Posit32::EncodeRegimeBits(Int32).0._State_7\;
                        end if;
                        
                    when \Posit32::EncodeRegimeBits(Int32).0._State_7\ => 
                        
                        \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.6\ := shift_left(\Posit32::EncodeRegimeBits(Int32).0.num\, to_integer(unsigned(SmartResize(\Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.5\, 5))));
                        \Posit32::EncodeRegimeBits(Int32).0.return\ <= \Posit32::EncodeRegimeBits(Int32).0.binaryOperationResult.6\;
                        \Posit32::EncodeRegimeBits(Int32).0._State\ := \Posit32::EncodeRegimeBits(Int32).0._State_1\;
                        
                        if (\Posit32::EncodeRegimeBits(Int32).0._State\ = \Posit32::EncodeRegimeBits(Int32).0._State_7\) then 
                            \Posit32::EncodeRegimeBits(Int32).0._State\ := \Posit32::EncodeRegimeBits(Int32).0._State_3\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._StateMachine\: process (\Clock\) 
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\: \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._States\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_0\;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.signBit\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.regimeKValue\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.1\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional080c1e8270378fd06e215f3c8f2add99c4865c1fbe8dd647a36c0c7e2edafab9\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.1\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.4\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.5\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional8ec324176b3f3fcd58fd5cfa6806fcab9222414090d26d94c66a65f1e77ad791\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.6\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.7\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.8\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.9\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.10\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.11\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalc44e6e18dba54d497a9ebfd5cd45c62d920ed273ec5aec35f89d9d27a8e797d3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalfaf425f73af9abdd07507acc85c797211aab0cbc36083f9065056c957f27c6b3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.12\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.13\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.14\: signed(63 downto 0) := to_signed(0, 64);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.15\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalb43e86d5d828dd5119f9f88af0ba7c790398b5cca8ee395bf1a45e5780b616e0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num3\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.4\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.16\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.5\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num4\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.17\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.18\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalbf654792f1ef201c91607ce88a255151da71234b0142c97b5e2a3594fec8b3f2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.19\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.20\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.21\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.22\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.23\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional0557e32b11ba8656de63af77389f74397db38458b6838b7ec71d9300b43b97b3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.24\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.25\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.26\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.27\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.28\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.29\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.30\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional18df916b486c957f6d73b71f963f462865051a4dad21055f9f7bb67a1b272e87\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.31\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.32\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.33\: signed(63 downto 0) := to_signed(0, 64);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.34\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionala777843480080cfd7ce563a33d79f12dd3aff5a7f1e7ee2bc6ae68dce3ba9f02\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.6\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._Finished\ <= false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return\ <= to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::EncodeRegimeBits(Int32).regimeKValue.parameter.Out.0\ <= to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::EncodeRegimeBits(Int32)._Started.0\ <= false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte).bits.parameter.Out.0\ <= to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte).startingPosition.parameter.Out.0\ <= to_unsigned(0, 8);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\ <= false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32).bits.parameter.Out.0\ <= to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32)._Started.0\ <= false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetMostSignificantOnePosition(UInt32).bits.parameter.Out.0\ <= to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Started.0\ <= false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::SetZero(UInt32,UInt16).bits.parameter.Out.0\ <= to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::SetZero(UInt32,UInt16).index.parameter.Out.0\ <= to_unsigned(0, 16);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::SetZero(UInt32,UInt16)._Started.0\ <= false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_0\;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.signBit\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.regimeKValue\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.0\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b\ := to_unsigned(0, 8);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.1\ := to_unsigned(0, 8);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.0\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional080c1e8270378fd06e215f3c8f2add99c4865c1fbe8dd647a36c0c7e2edafab9\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.1\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.2\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.0\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.3\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.4\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.5\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional8ec324176b3f3fcd58fd5cfa6806fcab9222414090d26d94c66a65f1e77ad791\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.6\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.7\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.8\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.9\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.10\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.11\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalc44e6e18dba54d497a9ebfd5cd45c62d920ed273ec5aec35f89d9d27a8e797d3\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.2\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalfaf425f73af9abdd07507acc85c797211aab0cbc36083f9065056c957f27c6b3\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.12\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.13\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.14\ := to_signed(0, 64);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.15\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalb43e86d5d828dd5119f9f88af0ba7c790398b5cca8ee395bf1a45e5780b616e0\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.3\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num3\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.4\ := to_unsigned(0, 8);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.16\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.5\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num4\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.17\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.18\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalbf654792f1ef201c91607ce88a255151da71234b0142c97b5e2a3594fec8b3f2\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.19\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.20\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.1\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.21\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.22\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.23\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional0557e32b11ba8656de63af77389f74397db38458b6838b7ec71d9300b43b97b3\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.24\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.25\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.26\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.2\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.27\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.28\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.29\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.30\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional18df916b486c957f6d73b71f963f462865051a4dad21055f9f7bb67a1b272e87\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.31\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.32\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.33\ := to_signed(0, 64);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.34\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionala777843480080cfd7ce563a33d79f12dd3aff5a7f1e7ee2bc6ae68dce3ba9f02\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.6\ := to_unsigned(0, 32);
            else 
                case \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ is 
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_0\ => 
                        
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._Started\ = true) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_2\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_1\ => 
                        
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._Started\ = true) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._Finished\ <= true;
                        else 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._Finished\ <= false;
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_0\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_2\ => 
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.signBit\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.signBit.parameter.In\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.regimeKValue\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.regimeKValue.parameter.In\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits.parameter.In\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits.parameter.In\;
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::EncodeRegimeBits(Int32).regimeKValue.parameter.Out.0\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.regimeKValue\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::EncodeRegimeBits(Int32)._Started.0\ <= true;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_3\;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_3\ => 
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::EncodeRegimeBits(Int32)._Started.0\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::EncodeRegimeBits(Int32)._Finished.0\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::EncodeRegimeBits(Int32)._Started.0\ <= false;
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.0\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::EncodeRegimeBits(Int32).return.0\;
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.0\;
                            
                            
                            
                            
                            
                            
                            
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte).bits.parameter.Out.0\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\;
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte).startingPosition.parameter.Out.0\ <= SmartResize(unsigned(to_signed(31, 32)), 8);
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\ <= true;
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_4\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_4\ => 
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\ <= false;
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.1\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte).return.0\;
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.1\;
                            
                            
                            
                            
                            
                            
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.0\ := to_signed(28, 32) - signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b\), 32));
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.0\);
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.1\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2\ >= to_signed(0, 32);

                            
                            
                            
                            

                            if ((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.1\)) then 
                                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_6\;
                            else 
                                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_7\;
                            end if;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_5\ => 
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.4\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\ + (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional080c1e8270378fd06e215f3c8f2add99c4865c1fbe8dd647a36c0c7e2edafab9\);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.4\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.5\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2\ < to_signed(0, 32);

                        
                        
                        

                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.5\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_9\;
                        else 
                            
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_8\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_6\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.2\ := shift_left(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits\, to_integer(unsigned(SmartResize(unsigned(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2\), 5))));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional080c1e8270378fd06e215f3c8f2add99c4865c1fbe8dd647a36c0c7e2edafab9\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.2\);
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_6\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_5\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_7\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.0\ := -\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.3\ := shift_right(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits\, to_integer(unsigned(SmartResize(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.0\, 5) and "11111")));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional080c1e8270378fd06e215f3c8f2add99c4865c1fbe8dd647a36c0c7e2edafab9\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.3\);
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_7\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_5\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_8\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetMostSignificantOnePosition(UInt32).bits.parameter.Out.0\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Started.0\ <= true;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_27\;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_9\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.6\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2\ > to_signed(28, 32);

                        
                        
                        
                        

                        if ((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.6\)) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_11\;
                        else 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_13\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_10\ => 
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional8ec324176b3f3fcd58fd5cfa6806fcab9222414090d26d94c66a65f1e77ad791\);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.11\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits\ < "10000000000000000000000000000000";

                        
                        
                        

                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.11\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_15\;
                        else 
                            
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_14\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_11\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.7\ := to_signed(32, 32) + \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_12\;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_12\ => 
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.8\ := shift_right(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits\, to_integer(unsigned(SmartResize(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.7\, 5) and "11111")));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional8ec324176b3f3fcd58fd5cfa6806fcab9222414090d26d94c66a65f1e77ad791\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.8\);
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_12\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_10\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_13\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.9\ := to_signed(32, 32) + \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.10\ := shift_left(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits\, to_integer(unsigned(SmartResize(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.9\, 5))));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional8ec324176b3f3fcd58fd5cfa6806fcab9222414090d26d94c66a65f1e77ad791\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.10\);
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_13\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_10\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_14\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.12\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits\ /= "10000000000000000000000000000000";

                        
                        
                        
                        

                        if ((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.12\)) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_21\;
                        else 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_22\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_15\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        

                        
                        
                        
                        

                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.signBit\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_17\;
                        else 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_19\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_16\ => 
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalc44e6e18dba54d497a9ebfd5cd45c62d920ed273ec5aec35f89d9d27a8e797d3\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_1\;
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_16\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_14\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_17\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32).bits.parameter.Out.0\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32)._Started.0\ <= true;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_18\;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_18\ => 
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32)._Started.0\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32)._Finished.0\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32)._Started.0\ <= false;
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.2\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32).return.0\;
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalc44e6e18dba54d497a9ebfd5cd45c62d920ed273ec5aec35f89d9d27a8e797d3\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.2\;
                            
                            if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_18\) then 
                                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_16\;
                            end if;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_19\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalc44e6e18dba54d497a9ebfd5cd45c62d920ed273ec5aec35f89d9d27a8e797d3\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\;
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_19\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_16\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_20\ => 
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalfaf425f73af9abdd07507acc85c797211aab0cbc36083f9065056c957f27c6b3\);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        

                        
                        
                        
                        

                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.signBit\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_24\;
                        else 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_26\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_21\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.13\ := SmartResize(unsigned(signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\), 64)) + to_signed(1, 64)), 32);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalfaf425f73af9abdd07507acc85c797211aab0cbc36083f9065056c957f27c6b3\ := ((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.13\));
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_21\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_20\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_22\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.14\ := signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\), 64)) and to_signed(1, 64);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.15\ := SmartResize(unsigned(signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\), 64)) + (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.14\)), 32);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalfaf425f73af9abdd07507acc85c797211aab0cbc36083f9065056c957f27c6b3\ := ((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.15\));
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_22\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_20\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_23\ => 
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalb43e86d5d828dd5119f9f88af0ba7c790398b5cca8ee395bf1a45e5780b616e0\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_1\;
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_23\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_8\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_24\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32).bits.parameter.Out.0\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32)._Started.0\ <= true;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_25\;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_25\ => 
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32)._Started.0\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32)._Finished.0\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32)._Started.0\ <= false;
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.3\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32).return.0\;
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalb43e86d5d828dd5119f9f88af0ba7c790398b5cca8ee395bf1a45e5780b616e0\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.3\;
                            
                            if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_25\) then 
                                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_23\;
                            end if;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_26\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalb43e86d5d828dd5119f9f88af0ba7c790398b5cca8ee395bf1a45e5780b616e0\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\;
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_26\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_23\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_27\ => 
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Started.0\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Finished.0\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Started.0\ <= false;
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.4\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetMostSignificantOnePosition(UInt32).return.0\;
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.16\ := signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.4\), 32)) - to_signed(1, 32);
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num3\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.16\);
                            
                            
                            
                            
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::SetZero(UInt32,UInt16).bits.parameter.Out.0\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\;
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::SetZero(UInt32,UInt16).index.parameter.Out.0\ <= SmartResize(unsigned(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num3\), 16);
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::SetZero(UInt32,UInt16)._Started.0\ <= true;
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_28\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_28\ => 
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::SetZero(UInt32,UInt16)._Started.0\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::SetZero(UInt32,UInt16)._Finished.0\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::SetZero(UInt32,UInt16)._Started.0\ <= false;
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.5\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::SetZero(UInt32,UInt16).return.0\;
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.5\;
                            
                            
                            
                            
                            
                            
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.17\ := to_signed(28, 32) - \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num3\;
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.18\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.17\) - signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b\), 32));
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num4\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.18\);
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_29\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_29\ => 
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.19\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num4\ >= to_signed(0, 32);

                        
                        
                        
                        

                        if ((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.19\)) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_31\;
                        else 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_32\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_30\ => 
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.22\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\ + (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalbf654792f1ef201c91607ce88a255151da71234b0142c97b5e2a3594fec8b3f2\);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.22\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.23\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num4\ < to_signed(0, 32);

                        
                        
                        

                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.23\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_34\;
                        else 
                            
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_33\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_31\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.20\ := shift_left(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\, to_integer(unsigned(SmartResize(unsigned(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num4\), 5))));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalbf654792f1ef201c91607ce88a255151da71234b0142c97b5e2a3594fec8b3f2\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.20\);
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_31\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_30\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_32\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.1\ := -\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num4\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.21\ := shift_right(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\, to_integer(unsigned(SmartResize(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.1\, 5) and "11111")));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalbf654792f1ef201c91607ce88a255151da71234b0142c97b5e2a3594fec8b3f2\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.21\);
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_32\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_30\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_33\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        

                        
                        
                        
                        

                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.signBit\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_45\;
                        else 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_47\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_34\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.24\ := to_signed(32, 32) + \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num4\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.25\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.24\ < to_signed(0, 32);

                        
                        
                        
                        

                        if ((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.25\)) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_36\;
                        else 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_38\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_35\ => 
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional0557e32b11ba8656de63af77389f74397db38458b6838b7ec71d9300b43b97b3\);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.30\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\ >= "10000000000000000000000000000000";

                        
                        
                        

                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.30\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_40\;
                        else 
                            
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_39\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_36\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.26\ := to_signed(32, 32) - \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num4\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.2\ := -(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.26\);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_37\;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_37\ => 
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.27\ := shift_right(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\, to_integer(unsigned(SmartResize(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.2\, 5) and "11111")));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional0557e32b11ba8656de63af77389f74397db38458b6838b7ec71d9300b43b97b3\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.27\);
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_37\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_35\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_38\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.28\ := to_signed(32, 32) + \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num4\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.29\ := shift_left(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\, to_integer(unsigned(SmartResize(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.28\, 5))));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional0557e32b11ba8656de63af77389f74397db38458b6838b7ec71d9300b43b97b3\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.29\);
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_38\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_35\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_39\ => 
                        
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_39\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_33\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_40\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.31\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\ /= "10000000000000000000000000000000";

                        
                        
                        
                        

                        if ((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.31\)) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_42\;
                        else 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_43\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_41\ => 
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional18df916b486c957f6d73b71f963f462865051a4dad21055f9f7bb67a1b272e87\);
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_41\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_39\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_42\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.32\ := SmartResize(unsigned(signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\), 64)) + to_signed(1, 64)), 32);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional18df916b486c957f6d73b71f963f462865051a4dad21055f9f7bb67a1b272e87\ := ((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.32\));
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_42\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_41\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_43\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.33\ := signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\), 64)) and to_signed(1, 64);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.34\ := SmartResize(unsigned(signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\), 64)) + (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.33\)), 32);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional18df916b486c957f6d73b71f963f462865051a4dad21055f9f7bb67a1b272e87\ := ((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.34\));
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_43\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_41\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_44\ => 
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionala777843480080cfd7ce563a33d79f12dd3aff5a7f1e7ee2bc6ae68dce3ba9f02\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_1\;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_45\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32).bits.parameter.Out.0\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32)._Started.0\ <= true;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_46\;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_46\ => 
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32)._Started.0\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32)._Finished.0\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32)._Started.0\ <= false;
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.6\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32).return.0\;
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionala777843480080cfd7ce563a33d79f12dd3aff5a7f1e7ee2bc6ae68dce3ba9f02\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return.6\;
                            
                            if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_46\) then 
                                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_44\;
                            end if;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_47\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionala777843480080cfd7ce563a33d79f12dd3aff5a7f1e7ee2bc6ae68dce3ba9f02\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\;
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_47\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_44\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::GetRegimeKValue().0._StateMachine\: process (\Clock\) 
        Variable \Posit32::GetRegimeKValue().0._State\: \Posit32::GetRegimeKValue().0._States\ := \Posit32::GetRegimeKValue().0._State_0\;
        Variable \Posit32::GetRegimeKValue().0.this\: \Lombiq.Arithmetics.Posit32\;
        Variable \Posit32::GetRegimeKValue().0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::GetRegimeKValue().0.conditional054ffdc2634715c514e630840f155e53d1c8ffe0be53ec06d4c21ba08ad2b716\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::GetRegimeKValue().0.b\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::GetRegimeKValue().0.return.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::GetRegimeKValue().0.conditional882cd98d817375e03765080fbf2e91fcc69740961af08057feb5bee6e57e0737\: signed(7 downto 0) := to_signed(0, 8);
        Variable \Posit32::GetRegimeKValue().0.unaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::GetRegimeKValue().0._Finished\ <= false;
                \Posit32::GetRegimeKValue().0.return\ <= to_signed(0, 8);
                \Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte).bits.parameter.Out.0\ <= to_unsigned(0, 32);
                \Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte).startingPosition.parameter.Out.0\ <= to_unsigned(0, 8);
                \Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\ <= false;
                \Posit32::GetRegimeKValue().0._State\ := \Posit32::GetRegimeKValue().0._State_0\;
                \Posit32::GetRegimeKValue().0.num\ := to_unsigned(0, 32);
                \Posit32::GetRegimeKValue().0.conditional054ffdc2634715c514e630840f155e53d1c8ffe0be53ec06d4c21ba08ad2b716\ := to_unsigned(0, 32);
                \Posit32::GetRegimeKValue().0.b\ := to_unsigned(0, 8);
                \Posit32::GetRegimeKValue().0.return.0\ := to_unsigned(0, 8);
                \Posit32::GetRegimeKValue().0.conditional882cd98d817375e03765080fbf2e91fcc69740961af08057feb5bee6e57e0737\ := to_signed(0, 8);
                \Posit32::GetRegimeKValue().0.unaryOperationResult.0\ := to_signed(0, 32);
            else 
                case \Posit32::GetRegimeKValue().0._State\ is 
                    when \Posit32::GetRegimeKValue().0._State_0\ => 
                        
                        
                        if (\Posit32::GetRegimeKValue().0._Started\ = true) then 
                            \Posit32::GetRegimeKValue().0._State\ := \Posit32::GetRegimeKValue().0._State_2\;
                        end if;
                        
                    when \Posit32::GetRegimeKValue().0._State_1\ => 
                        
                        
                        if (\Posit32::GetRegimeKValue().0._Started\ = true) then 
                            \Posit32::GetRegimeKValue().0._Finished\ <= true;
                        else 
                            \Posit32::GetRegimeKValue().0._Finished\ <= false;
                            \Posit32::GetRegimeKValue().0._State\ := \Posit32::GetRegimeKValue().0._State_0\;
                        end if;
                        
                    when \Posit32::GetRegimeKValue().0._State_2\ => 
                        \Posit32::GetRegimeKValue().0.this\ := \Posit32::GetRegimeKValue().0.this.parameter.In\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::GetRegimeKValue().0.conditional054ffdc2634715c514e630840f155e53d1c8ffe0be53ec06d4c21ba08ad2b716\ := to_unsigned(0, 32);
                        
                        
                        
                        \Posit32::GetRegimeKValue().0.num\ := to_unsigned(0, 32);
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte).bits.parameter.Out.0\ <= to_unsigned(0, 32);
                        \Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte).startingPosition.parameter.Out.0\ <= SmartResize(unsigned(to_signed(31, 32)), 8);
                        \Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\ <= true;
                        \Posit32::GetRegimeKValue().0._State\ := \Posit32::GetRegimeKValue().0._State_3\;
                        
                    when \Posit32::GetRegimeKValue().0._State_3\ => 
                        
                        if (\Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\ = \Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\) then 
                            \Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\ <= false;
                            \Posit32::GetRegimeKValue().0.return.0\ := \Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte).return.0\;
                            \Posit32::GetRegimeKValue().0.b\ := \Posit32::GetRegimeKValue().0.return.0\;
                            
                            
                            
                            
                            
                            
                            \Posit32::GetRegimeKValue().0.unaryOperationResult.0\ := -signed(SmartResize((\Posit32::GetRegimeKValue().0.b\), 32));
                            \Posit32::GetRegimeKValue().0.conditional882cd98d817375e03765080fbf2e91fcc69740961af08057feb5bee6e57e0737\ := (SmartResize((\Posit32::GetRegimeKValue().0.unaryOperationResult.0\), 8));
                            
                            
                            
                            \Posit32::GetRegimeKValue().0.return\ <= \Posit32::GetRegimeKValue().0.conditional882cd98d817375e03765080fbf2e91fcc69740961af08057feb5bee6e57e0737\;
                            \Posit32::GetRegimeKValue().0._State\ := \Posit32::GetRegimeKValue().0._State_1\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::CalculateScaleFactor().0._StateMachine\: process (\Clock\) 
        Variable \Posit32::CalculateScaleFactor().0._State\: \Posit32::CalculateScaleFactor().0._States\ := \Posit32::CalculateScaleFactor().0._State_0\;
        Variable \Posit32::CalculateScaleFactor().0.this\: \Lombiq.Arithmetics.Posit32\;
        Variable \Posit32::CalculateScaleFactor().0.regimeKValue\: signed(7 downto 0) := to_signed(0, 8);
        Variable \Posit32::CalculateScaleFactor().0.return.0\: signed(7 downto 0) := to_signed(0, 8);
        Variable \Posit32::CalculateScaleFactor().0.conditional1aa95b35288eb627929161a1ee637479589960934567100c958634e64afb13de\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::CalculateScaleFactor().0.binaryOperationResult.0\: boolean := false;
        Variable \Posit32::CalculateScaleFactor().0.binaryOperationResult.1\: signed(63 downto 0) := to_signed(0, 64);
        Variable \Posit32::CalculateScaleFactor().0.return.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::CalculateScaleFactor().0.binaryOperationResult.2\: signed(15 downto 0) := to_signed(0, 16);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::CalculateScaleFactor().0._Finished\ <= false;
                \Posit32::CalculateScaleFactor().0.return\ <= to_signed(0, 16);
                \Posit32::CalculateScaleFactor().0.Posit32::GetRegimeKValue()._Started.0\ <= false;
                \Posit32::CalculateScaleFactor().0.Posit32::GetExponentValue()._Started.0\ <= false;
                \Posit32::CalculateScaleFactor().0._State\ := \Posit32::CalculateScaleFactor().0._State_0\;
                \Posit32::CalculateScaleFactor().0.regimeKValue\ := to_signed(0, 8);
                \Posit32::CalculateScaleFactor().0.return.0\ := to_signed(0, 8);
                \Posit32::CalculateScaleFactor().0.conditional1aa95b35288eb627929161a1ee637479589960934567100c958634e64afb13de\ := to_signed(0, 32);
                \Posit32::CalculateScaleFactor().0.binaryOperationResult.0\ := false;
                \Posit32::CalculateScaleFactor().0.binaryOperationResult.1\ := to_signed(0, 64);
                \Posit32::CalculateScaleFactor().0.return.1\ := to_unsigned(0, 32);
                \Posit32::CalculateScaleFactor().0.binaryOperationResult.2\ := to_signed(0, 16);
            else 
                case \Posit32::CalculateScaleFactor().0._State\ is 
                    when \Posit32::CalculateScaleFactor().0._State_0\ => 
                        
                        
                        if (\Posit32::CalculateScaleFactor().0._Started\ = true) then 
                            \Posit32::CalculateScaleFactor().0._State\ := \Posit32::CalculateScaleFactor().0._State_2\;
                        end if;
                        
                    when \Posit32::CalculateScaleFactor().0._State_1\ => 
                        
                        
                        if (\Posit32::CalculateScaleFactor().0._Started\ = true) then 
                            \Posit32::CalculateScaleFactor().0._Finished\ <= true;
                        else 
                            \Posit32::CalculateScaleFactor().0._Finished\ <= false;
                            \Posit32::CalculateScaleFactor().0._State\ := \Posit32::CalculateScaleFactor().0._State_0\;
                        end if;
                        
                    when \Posit32::CalculateScaleFactor().0._State_2\ => 
                        \Posit32::CalculateScaleFactor().0.this\ := \Posit32::CalculateScaleFactor().0.this.parameter.In\;
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::CalculateScaleFactor().0.Posit32::GetRegimeKValue().this.parameter.Out.0\ <= \Posit32::CalculateScaleFactor().0.this\;
                        \Posit32::CalculateScaleFactor().0.Posit32::GetRegimeKValue()._Started.0\ <= true;
                        \Posit32::CalculateScaleFactor().0._State\ := \Posit32::CalculateScaleFactor().0._State_3\;
                        
                    when \Posit32::CalculateScaleFactor().0._State_3\ => 
                        
                        if (\Posit32::CalculateScaleFactor().0.Posit32::GetRegimeKValue()._Started.0\ = \Posit32::CalculateScaleFactor().0.Posit32::GetRegimeKValue()._Finished.0\) then 
                            \Posit32::CalculateScaleFactor().0.Posit32::GetRegimeKValue()._Started.0\ <= false;
                            \Posit32::CalculateScaleFactor().0.return.0\ := \Posit32::CalculateScaleFactor().0.Posit32::GetRegimeKValue().return.0\;
                            \Posit32::CalculateScaleFactor().0.regimeKValue\ := \Posit32::CalculateScaleFactor().0.return.0\;
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32::CalculateScaleFactor().0.binaryOperationResult.0\ := SmartResize((\Posit32::CalculateScaleFactor().0.regimeKValue\), 32) /= to_signed(-31, 32);

                            
                            
                            
                            

                            if ((\Posit32::CalculateScaleFactor().0.binaryOperationResult.0\)) then 
                                \Posit32::CalculateScaleFactor().0._State\ := \Posit32::CalculateScaleFactor().0._State_5\;
                            else 
                                \Posit32::CalculateScaleFactor().0._State\ := \Posit32::CalculateScaleFactor().0._State_7\;
                            end if;
                        end if;
                        
                    when \Posit32::CalculateScaleFactor().0._State_4\ => 
                        
                        
                        
                        
                        \Posit32::CalculateScaleFactor().0.return\ <= SmartResize((\Posit32::CalculateScaleFactor().0.conditional1aa95b35288eb627929161a1ee637479589960934567100c958634e64afb13de\), 16);
                        \Posit32::CalculateScaleFactor().0._State\ := \Posit32::CalculateScaleFactor().0._State_1\;
                        
                    when \Posit32::CalculateScaleFactor().0._State_5\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::CalculateScaleFactor().0.binaryOperationResult.1\ := SmartResize(SmartResize((\Posit32::CalculateScaleFactor().0.regimeKValue\), 32) * to_signed(4, 32), 64);
                        
                        \Posit32::CalculateScaleFactor().0.Posit32::GetExponentValue().this.parameter.Out.0\ <= \Posit32::CalculateScaleFactor().0.this\;
                        \Posit32::CalculateScaleFactor().0.Posit32::GetExponentValue()._Started.0\ <= true;
                        \Posit32::CalculateScaleFactor().0._State\ := \Posit32::CalculateScaleFactor().0._State_6\;
                        
                    when \Posit32::CalculateScaleFactor().0._State_6\ => 
                        
                        if (\Posit32::CalculateScaleFactor().0.Posit32::GetExponentValue()._Started.0\ = \Posit32::CalculateScaleFactor().0.Posit32::GetExponentValue()._Finished.0\) then 
                            \Posit32::CalculateScaleFactor().0.Posit32::GetExponentValue()._Started.0\ <= false;
                            \Posit32::CalculateScaleFactor().0.return.1\ := \Posit32::CalculateScaleFactor().0.Posit32::GetExponentValue().return.0\;
                            \Posit32::CalculateScaleFactor().0.binaryOperationResult.2\ := SmartResize((\Posit32::CalculateScaleFactor().0.binaryOperationResult.1\) + signed(SmartResize((\Posit32::CalculateScaleFactor().0.return.1\), 64)), 16);
                            \Posit32::CalculateScaleFactor().0.conditional1aa95b35288eb627929161a1ee637479589960934567100c958634e64afb13de\ := SmartResize(((\Posit32::CalculateScaleFactor().0.binaryOperationResult.2\)), 32);
                            
                            if (\Posit32::CalculateScaleFactor().0._State\ = \Posit32::CalculateScaleFactor().0._State_6\) then 
                                \Posit32::CalculateScaleFactor().0._State\ := \Posit32::CalculateScaleFactor().0._State_4\;
                            end if;
                        end if;
                        
                    when \Posit32::CalculateScaleFactor().0._State_7\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::CalculateScaleFactor().0.conditional1aa95b35288eb627929161a1ee637479589960934567100c958634e64afb13de\ := to_signed(0, 32);
                        
                        if (\Posit32::CalculateScaleFactor().0._State\ = \Posit32::CalculateScaleFactor().0._State_7\) then 
                            \Posit32::CalculateScaleFactor().0._State\ := \Posit32::CalculateScaleFactor().0._State_4\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::ExponentSize().0._StateMachine\: process (\Clock\) 
        Variable \Posit32::ExponentSize().0._State\: \Posit32::ExponentSize().0._States\ := \Posit32::ExponentSize().0._State_0\;
        Variable \Posit32::ExponentSize().0.this\: \Lombiq.Arithmetics.Posit32\;
        Variable \Posit32::ExponentSize().0.bits\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::ExponentSize().0.conditional85ca8d8893aa24483d9e74ed87417b722b6d33d6069def85ee5195c77759eab3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::ExponentSize().0.b\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::ExponentSize().0.return.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::ExponentSize().0.binaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::ExponentSize().0.binaryOperationResult.1\: boolean := false;
        Variable \Posit32::ExponentSize().0.conditional68bcd4673000ed90d5e5bddf9742548ff8843dd36c272b449a1de261af0ae5a9\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::ExponentSize().0.binaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::ExponentSize().0.binaryOperationResult.3\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::ExponentSize().0.binaryOperationResult.4\: boolean := false;
        Variable \Posit32::ExponentSize().0.binaryOperationResult.5\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::ExponentSize().0.binaryOperationResult.6\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::ExponentSize().0.binaryOperationResult.7\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::ExponentSize().0.binaryOperationResult.8\: unsigned(7 downto 0) := to_unsigned(0, 8);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::ExponentSize().0._Finished\ <= false;
                \Posit32::ExponentSize().0.return\ <= to_unsigned(0, 8);
                \Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte).bits.parameter.Out.0\ <= to_unsigned(0, 32);
                \Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte).startingPosition.parameter.Out.0\ <= to_unsigned(0, 8);
                \Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\ <= false;
                \Posit32::ExponentSize().0._State\ := \Posit32::ExponentSize().0._State_0\;
                \Posit32::ExponentSize().0.bits\ := to_unsigned(0, 32);
                \Posit32::ExponentSize().0.conditional85ca8d8893aa24483d9e74ed87417b722b6d33d6069def85ee5195c77759eab3\ := to_unsigned(0, 32);
                \Posit32::ExponentSize().0.b\ := to_unsigned(0, 8);
                \Posit32::ExponentSize().0.return.0\ := to_unsigned(0, 8);
                \Posit32::ExponentSize().0.binaryOperationResult.0\ := to_signed(0, 32);
                \Posit32::ExponentSize().0.binaryOperationResult.1\ := false;
                \Posit32::ExponentSize().0.conditional68bcd4673000ed90d5e5bddf9742548ff8843dd36c272b449a1de261af0ae5a9\ := to_signed(0, 32);
                \Posit32::ExponentSize().0.binaryOperationResult.2\ := to_signed(0, 32);
                \Posit32::ExponentSize().0.binaryOperationResult.3\ := to_signed(0, 32);
                \Posit32::ExponentSize().0.binaryOperationResult.4\ := false;
                \Posit32::ExponentSize().0.binaryOperationResult.5\ := to_signed(0, 32);
                \Posit32::ExponentSize().0.binaryOperationResult.6\ := to_unsigned(0, 8);
                \Posit32::ExponentSize().0.binaryOperationResult.7\ := to_signed(0, 32);
                \Posit32::ExponentSize().0.binaryOperationResult.8\ := to_unsigned(0, 8);
            else 
                case \Posit32::ExponentSize().0._State\ is 
                    when \Posit32::ExponentSize().0._State_0\ => 
                        
                        
                        if (\Posit32::ExponentSize().0._Started\ = true) then 
                            \Posit32::ExponentSize().0._State\ := \Posit32::ExponentSize().0._State_2\;
                        end if;
                        
                    when \Posit32::ExponentSize().0._State_1\ => 
                        
                        
                        if (\Posit32::ExponentSize().0._Started\ = true) then 
                            \Posit32::ExponentSize().0._Finished\ <= true;
                        else 
                            \Posit32::ExponentSize().0._Finished\ <= false;
                            \Posit32::ExponentSize().0._State\ := \Posit32::ExponentSize().0._State_0\;
                        end if;
                        
                    when \Posit32::ExponentSize().0._State_2\ => 
                        \Posit32::ExponentSize().0.this\ := \Posit32::ExponentSize().0.this.parameter.In\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::ExponentSize().0.conditional85ca8d8893aa24483d9e74ed87417b722b6d33d6069def85ee5195c77759eab3\ := to_unsigned(0, 32);
                        
                        
                        
                        \Posit32::ExponentSize().0.bits\ := to_unsigned(0, 32);
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte).bits.parameter.Out.0\ <= to_unsigned(0, 32);
                        \Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte).startingPosition.parameter.Out.0\ <= SmartResize(unsigned(to_signed(31, 32)), 8);
                        \Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\ <= true;
                        \Posit32::ExponentSize().0._State\ := \Posit32::ExponentSize().0._State_3\;
                        
                    when \Posit32::ExponentSize().0._State_3\ => 
                        
                        if (\Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\ = \Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\) then 
                            \Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\ <= false;
                            \Posit32::ExponentSize().0.return.0\ := \Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte).return.0\;
                            \Posit32::ExponentSize().0.b\ := \Posit32::ExponentSize().0.return.0\;
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32::ExponentSize().0.binaryOperationResult.0\ := signed(SmartResize((\Posit32::ExponentSize().0.b\), 32)) + to_signed(2, 32);
                            \Posit32::ExponentSize().0.binaryOperationResult.1\ := \Posit32::ExponentSize().0.binaryOperationResult.0\ <= to_signed(32, 32);

                            
                            
                            

                            if (\Posit32::ExponentSize().0.binaryOperationResult.1\) then 
                                \Posit32::ExponentSize().0._State\ := \Posit32::ExponentSize().0._State_5\;
                            else 
                                
                                \Posit32::ExponentSize().0._State\ := \Posit32::ExponentSize().0._State_4\;
                            end if;
                        end if;
                        
                    when \Posit32::ExponentSize().0._State_4\ => 
                        
                        
                        
                        
                        \Posit32::ExponentSize().0.binaryOperationResult.7\ := to_signed(32, 32) - signed(SmartResize((\Posit32::ExponentSize().0.b\), 32));
                        \Posit32::ExponentSize().0.binaryOperationResult.8\ := SmartResize(unsigned(\Posit32::ExponentSize().0.binaryOperationResult.7\ - to_signed(1, 32)), 8);
                        \Posit32::ExponentSize().0.return\ <= (\Posit32::ExponentSize().0.binaryOperationResult.8\);
                        \Posit32::ExponentSize().0._State\ := \Posit32::ExponentSize().0._State_1\;
                        
                    when \Posit32::ExponentSize().0._State_5\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::ExponentSize().0.binaryOperationResult.2\ := signed(SmartResize((\Posit32::ExponentSize().0.b\), 32)) + to_signed(2, 32);
                        \Posit32::ExponentSize().0.binaryOperationResult.3\ := to_signed(32, 32) - (\Posit32::ExponentSize().0.binaryOperationResult.2\);
                        \Posit32::ExponentSize().0._State\ := \Posit32::ExponentSize().0._State_6\;
                        
                    when \Posit32::ExponentSize().0._State_6\ => 
                        
                        \Posit32::ExponentSize().0.binaryOperationResult.4\ := \Posit32::ExponentSize().0.binaryOperationResult.3\ > to_signed(2, 32);

                        
                        
                        
                        

                        if ((\Posit32::ExponentSize().0.binaryOperationResult.4\)) then 
                            \Posit32::ExponentSize().0._State\ := \Posit32::ExponentSize().0._State_8\;
                        else 
                            \Posit32::ExponentSize().0._State\ := \Posit32::ExponentSize().0._State_9\;
                        end if;
                        
                    when \Posit32::ExponentSize().0._State_7\ => 
                        
                        
                        
                        
                        \Posit32::ExponentSize().0.return\ <= SmartResize(unsigned((\Posit32::ExponentSize().0.conditional68bcd4673000ed90d5e5bddf9742548ff8843dd36c272b449a1de261af0ae5a9\)), 8);
                        \Posit32::ExponentSize().0._State\ := \Posit32::ExponentSize().0._State_1\;
                        
                        if (\Posit32::ExponentSize().0._State\ = \Posit32::ExponentSize().0._State_7\) then 
                            \Posit32::ExponentSize().0._State\ := \Posit32::ExponentSize().0._State_4\;
                        end if;
                        
                    when \Posit32::ExponentSize().0._State_8\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::ExponentSize().0.conditional68bcd4673000ed90d5e5bddf9742548ff8843dd36c272b449a1de261af0ae5a9\ := to_signed(2, 32);
                        
                        if (\Posit32::ExponentSize().0._State\ = \Posit32::ExponentSize().0._State_8\) then 
                            \Posit32::ExponentSize().0._State\ := \Posit32::ExponentSize().0._State_7\;
                        end if;
                        
                    when \Posit32::ExponentSize().0._State_9\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::ExponentSize().0.binaryOperationResult.5\ := signed(SmartResize((\Posit32::ExponentSize().0.b\), 32)) + to_signed(2, 32);
                        \Posit32::ExponentSize().0.binaryOperationResult.6\ := SmartResize(unsigned(to_signed(32, 32) - (\Posit32::ExponentSize().0.binaryOperationResult.5\)), 8);
                        \Posit32::ExponentSize().0.conditional68bcd4673000ed90d5e5bddf9742548ff8843dd36c272b449a1de261af0ae5a9\ := signed(SmartResize(((\Posit32::ExponentSize().0.binaryOperationResult.6\)), 32));
                        
                        if (\Posit32::ExponentSize().0._State\ = \Posit32::ExponentSize().0._State_9\) then 
                            \Posit32::ExponentSize().0._State\ := \Posit32::ExponentSize().0._State_7\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::GetExponentValue().0._StateMachine\: process (\Clock\) 
        Variable \Posit32::GetExponentValue().0._State\: \Posit32::GetExponentValue().0._States\ := \Posit32::GetExponentValue().0._State_0\;
        Variable \Posit32::GetExponentValue().0.this\: \Lombiq.Arithmetics.Posit32\;
        Variable \Posit32::GetExponentValue().0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::GetExponentValue().0.conditional880d0f3a8d33b2428fb4e8a62e4174f93b0cc01cc9b8d6d16563b7d2d4e90992\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::GetExponentValue().0.b\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::GetExponentValue().0.return.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::GetExponentValue().0.return.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::GetExponentValue().0.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::GetExponentValue().0.binaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::GetExponentValue().0.binaryOperationResult.2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::GetExponentValue().0.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::GetExponentValue().0.conditionala233560fe7dfff22c231bec46671f442fee11494dc774056e64d669ec36cdb00\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::GetExponentValue().0.binaryOperationResult.4\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::GetExponentValue().0._Finished\ <= false;
                \Posit32::GetExponentValue().0.return\ <= to_unsigned(0, 32);
                \Posit32::GetExponentValue().0.Posit32::ExponentSize()._Started.0\ <= false;
                \Posit32::GetExponentValue().0.Posit32::FractionSize()._Started.0\ <= false;
                \Posit32::GetExponentValue().0._State\ := \Posit32::GetExponentValue().0._State_0\;
                \Posit32::GetExponentValue().0.num\ := to_unsigned(0, 32);
                \Posit32::GetExponentValue().0.conditional880d0f3a8d33b2428fb4e8a62e4174f93b0cc01cc9b8d6d16563b7d2d4e90992\ := to_unsigned(0, 32);
                \Posit32::GetExponentValue().0.b\ := to_unsigned(0, 8);
                \Posit32::GetExponentValue().0.return.0\ := to_unsigned(0, 8);
                \Posit32::GetExponentValue().0.return.1\ := to_unsigned(0, 32);
                \Posit32::GetExponentValue().0.binaryOperationResult.0\ := to_unsigned(0, 32);
                \Posit32::GetExponentValue().0.binaryOperationResult.1\ := to_signed(0, 32);
                \Posit32::GetExponentValue().0.binaryOperationResult.2\ := to_unsigned(0, 32);
                \Posit32::GetExponentValue().0.binaryOperationResult.3\ := to_unsigned(0, 32);
                \Posit32::GetExponentValue().0.conditionala233560fe7dfff22c231bec46671f442fee11494dc774056e64d669ec36cdb00\ := to_unsigned(0, 32);
                \Posit32::GetExponentValue().0.binaryOperationResult.4\ := false;
            else 
                case \Posit32::GetExponentValue().0._State\ is 
                    when \Posit32::GetExponentValue().0._State_0\ => 
                        
                        
                        if (\Posit32::GetExponentValue().0._Started\ = true) then 
                            \Posit32::GetExponentValue().0._State\ := \Posit32::GetExponentValue().0._State_2\;
                        end if;
                        
                    when \Posit32::GetExponentValue().0._State_1\ => 
                        
                        
                        if (\Posit32::GetExponentValue().0._Started\ = true) then 
                            \Posit32::GetExponentValue().0._Finished\ <= true;
                        else 
                            \Posit32::GetExponentValue().0._Finished\ <= false;
                            \Posit32::GetExponentValue().0._State\ := \Posit32::GetExponentValue().0._State_0\;
                        end if;
                        
                    when \Posit32::GetExponentValue().0._State_2\ => 
                        \Posit32::GetExponentValue().0.this\ := \Posit32::GetExponentValue().0.this.parameter.In\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::GetExponentValue().0.conditional880d0f3a8d33b2428fb4e8a62e4174f93b0cc01cc9b8d6d16563b7d2d4e90992\ := to_unsigned(0, 32);
                        
                        
                        
                        \Posit32::GetExponentValue().0.num\ := to_unsigned(0, 32);
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::GetExponentValue().0.Posit32::ExponentSize().this.parameter.Out.0\ <= \Posit32::GetExponentValue().0.this\;
                        \Posit32::GetExponentValue().0.Posit32::ExponentSize()._Started.0\ <= true;
                        \Posit32::GetExponentValue().0._State\ := \Posit32::GetExponentValue().0._State_3\;
                        
                    when \Posit32::GetExponentValue().0._State_3\ => 
                        
                        if (\Posit32::GetExponentValue().0.Posit32::ExponentSize()._Started.0\ = \Posit32::GetExponentValue().0.Posit32::ExponentSize()._Finished.0\) then 
                            \Posit32::GetExponentValue().0.Posit32::ExponentSize()._Started.0\ <= false;
                            \Posit32::GetExponentValue().0.return.0\ := \Posit32::GetExponentValue().0.Posit32::ExponentSize().return.0\;
                            \Posit32::GetExponentValue().0.b\ := \Posit32::GetExponentValue().0.return.0\;
                            
                            
                            
                            
                            \Posit32::GetExponentValue().0.Posit32::FractionSize().this.parameter.Out.0\ <= \Posit32::GetExponentValue().0.this\;
                            \Posit32::GetExponentValue().0.Posit32::FractionSize()._Started.0\ <= true;
                            \Posit32::GetExponentValue().0._State\ := \Posit32::GetExponentValue().0._State_4\;
                        end if;
                        
                    when \Posit32::GetExponentValue().0._State_4\ => 
                        
                        if (\Posit32::GetExponentValue().0.Posit32::FractionSize()._Started.0\ = \Posit32::GetExponentValue().0.Posit32::FractionSize()._Finished.0\) then 
                            \Posit32::GetExponentValue().0.Posit32::FractionSize()._Started.0\ <= false;
                            \Posit32::GetExponentValue().0.return.1\ := \Posit32::GetExponentValue().0.Posit32::FractionSize().return.0\;
                            \Posit32::GetExponentValue().0.binaryOperationResult.0\ := shift_right(to_unsigned(0, 32), to_integer(unsigned(SmartResize(signed(\Posit32::GetExponentValue().0.return.1\), 5) and "11111")));
                            \Posit32::GetExponentValue().0.binaryOperationResult.1\ := to_signed(32, 32) - signed(SmartResize((\Posit32::GetExponentValue().0.b\), 32));
                            \Posit32::GetExponentValue().0._State\ := \Posit32::GetExponentValue().0._State_5\;
                        end if;
                        
                    when \Posit32::GetExponentValue().0._State_5\ => 
                        
                        \Posit32::GetExponentValue().0.binaryOperationResult.2\ := shift_left(\Posit32::GetExponentValue().0.binaryOperationResult.0\, to_integer(unsigned(SmartResize(\Posit32::GetExponentValue().0.binaryOperationResult.1\, 5))));
                        \Posit32::GetExponentValue().0.binaryOperationResult.3\ := shift_right(\Posit32::GetExponentValue().0.binaryOperationResult.2\, to_integer(unsigned(SmartResize(to_signed(30, 32), 5) and "11111")));
                        \Posit32::GetExponentValue().0.num\ := \Posit32::GetExponentValue().0.binaryOperationResult.3\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::GetExponentValue().0._State\ := \Posit32::GetExponentValue().0._State_6\;
                        
                    when \Posit32::GetExponentValue().0._State_6\ => 
                        
                        \Posit32::GetExponentValue().0.binaryOperationResult.4\ := signed(SmartResize((\Posit32::GetExponentValue().0.b\), 32)) /= to_signed(0, 32);

                        
                        
                        
                        

                        if ((\Posit32::GetExponentValue().0.binaryOperationResult.4\)) then 
                            \Posit32::GetExponentValue().0._State\ := \Posit32::GetExponentValue().0._State_8\;
                        else 
                            \Posit32::GetExponentValue().0._State\ := \Posit32::GetExponentValue().0._State_9\;
                        end if;
                        
                    when \Posit32::GetExponentValue().0._State_7\ => 
                        
                        
                        
                        
                        \Posit32::GetExponentValue().0.return\ <= \Posit32::GetExponentValue().0.conditionala233560fe7dfff22c231bec46671f442fee11494dc774056e64d669ec36cdb00\;
                        \Posit32::GetExponentValue().0._State\ := \Posit32::GetExponentValue().0._State_1\;
                        
                    when \Posit32::GetExponentValue().0._State_8\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::GetExponentValue().0.conditionala233560fe7dfff22c231bec46671f442fee11494dc774056e64d669ec36cdb00\ := \Posit32::GetExponentValue().0.num\;
                        
                        if (\Posit32::GetExponentValue().0._State\ = \Posit32::GetExponentValue().0._State_8\) then 
                            \Posit32::GetExponentValue().0._State\ := \Posit32::GetExponentValue().0._State_7\;
                        end if;
                        
                    when \Posit32::GetExponentValue().0._State_9\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::GetExponentValue().0.conditionala233560fe7dfff22c231bec46671f442fee11494dc774056e64d669ec36cdb00\ := to_unsigned(0, 32);
                        
                        if (\Posit32::GetExponentValue().0._State\ = \Posit32::GetExponentValue().0._State_9\) then 
                            \Posit32::GetExponentValue().0._State\ := \Posit32::GetExponentValue().0._State_7\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::FractionSize().0._StateMachine\: process (\Clock\) 
        Variable \Posit32::FractionSize().0._State\: \Posit32::FractionSize().0._States\ := \Posit32::FractionSize().0._State_0\;
        Variable \Posit32::FractionSize().0.this\: \Lombiq.Arithmetics.Posit32\;
        Variable \Posit32::FractionSize().0.bits\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::FractionSize().0.conditional963d17004b6788ad55358cce58986fa179ec1b5dc039dfede93d706448099e92\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::FractionSize().0.num\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::FractionSize().0.return.0\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::FractionSize().0.binaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::FractionSize().0.binaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::FractionSize().0.binaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::FractionSize().0.conditionalf2eba7c459dd057c9270f346c2a9013399b4309fc21683746ef1be47061f03f1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::FractionSize().0.binaryOperationResult.3\: boolean := false;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::FractionSize().0._Finished\ <= false;
                \Posit32::FractionSize().0.return\ <= to_unsigned(0, 32);
                \Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte).bits.parameter.Out.0\ <= to_unsigned(0, 32);
                \Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte).startingPosition.parameter.Out.0\ <= to_unsigned(0, 8);
                \Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\ <= false;
                \Posit32::FractionSize().0._State\ := \Posit32::FractionSize().0._State_0\;
                \Posit32::FractionSize().0.bits\ := to_unsigned(0, 32);
                \Posit32::FractionSize().0.conditional963d17004b6788ad55358cce58986fa179ec1b5dc039dfede93d706448099e92\ := to_unsigned(0, 32);
                \Posit32::FractionSize().0.num\ := to_signed(0, 32);
                \Posit32::FractionSize().0.return.0\ := to_unsigned(0, 8);
                \Posit32::FractionSize().0.binaryOperationResult.0\ := to_signed(0, 32);
                \Posit32::FractionSize().0.binaryOperationResult.1\ := to_signed(0, 32);
                \Posit32::FractionSize().0.binaryOperationResult.2\ := to_signed(0, 32);
                \Posit32::FractionSize().0.conditionalf2eba7c459dd057c9270f346c2a9013399b4309fc21683746ef1be47061f03f1\ := to_unsigned(0, 32);
                \Posit32::FractionSize().0.binaryOperationResult.3\ := false;
            else 
                case \Posit32::FractionSize().0._State\ is 
                    when \Posit32::FractionSize().0._State_0\ => 
                        
                        
                        if (\Posit32::FractionSize().0._Started\ = true) then 
                            \Posit32::FractionSize().0._State\ := \Posit32::FractionSize().0._State_2\;
                        end if;
                        
                    when \Posit32::FractionSize().0._State_1\ => 
                        
                        
                        if (\Posit32::FractionSize().0._Started\ = true) then 
                            \Posit32::FractionSize().0._Finished\ <= true;
                        else 
                            \Posit32::FractionSize().0._Finished\ <= false;
                            \Posit32::FractionSize().0._State\ := \Posit32::FractionSize().0._State_0\;
                        end if;
                        
                    when \Posit32::FractionSize().0._State_2\ => 
                        \Posit32::FractionSize().0.this\ := \Posit32::FractionSize().0.this.parameter.In\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::FractionSize().0.conditional963d17004b6788ad55358cce58986fa179ec1b5dc039dfede93d706448099e92\ := to_unsigned(0, 32);
                        
                        
                        
                        \Posit32::FractionSize().0.bits\ := to_unsigned(0, 32);
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte).bits.parameter.Out.0\ <= to_unsigned(0, 32);
                        \Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte).startingPosition.parameter.Out.0\ <= SmartResize(unsigned(to_signed(31, 32)), 8);
                        \Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\ <= true;
                        \Posit32::FractionSize().0._State\ := \Posit32::FractionSize().0._State_3\;
                        
                    when \Posit32::FractionSize().0._State_3\ => 
                        
                        if (\Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\ = \Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\) then 
                            \Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\ <= false;
                            \Posit32::FractionSize().0.return.0\ := \Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte).return.0\;
                            \Posit32::FractionSize().0.binaryOperationResult.0\ := signed(SmartResize((\Posit32::FractionSize().0.return.0\), 32)) + to_signed(2, 32);
                            \Posit32::FractionSize().0.binaryOperationResult.1\ := SmartResize(\Posit32::FractionSize().0.binaryOperationResult.0\ + to_signed(2, 32), 32);
                            \Posit32::FractionSize().0._State\ := \Posit32::FractionSize().0._State_4\;
                        end if;
                        
                    when \Posit32::FractionSize().0._State_4\ => 
                        
                        \Posit32::FractionSize().0.binaryOperationResult.2\ := to_signed(32, 32) - (\Posit32::FractionSize().0.binaryOperationResult.1\);
                        \Posit32::FractionSize().0.num\ := \Posit32::FractionSize().0.binaryOperationResult.2\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::FractionSize().0.binaryOperationResult.3\ := \Posit32::FractionSize().0.num\ > to_signed(0, 32);

                        
                        
                        
                        

                        if ((\Posit32::FractionSize().0.binaryOperationResult.3\)) then 
                            \Posit32::FractionSize().0._State\ := \Posit32::FractionSize().0._State_6\;
                        else 
                            \Posit32::FractionSize().0._State\ := \Posit32::FractionSize().0._State_7\;
                        end if;
                        
                    when \Posit32::FractionSize().0._State_5\ => 
                        
                        
                        
                        
                        \Posit32::FractionSize().0.return\ <= \Posit32::FractionSize().0.conditionalf2eba7c459dd057c9270f346c2a9013399b4309fc21683746ef1be47061f03f1\;
                        \Posit32::FractionSize().0._State\ := \Posit32::FractionSize().0._State_1\;
                        
                    when \Posit32::FractionSize().0._State_6\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::FractionSize().0.conditionalf2eba7c459dd057c9270f346c2a9013399b4309fc21683746ef1be47061f03f1\ := (unsigned(\Posit32::FractionSize().0.num\));
                        
                        if (\Posit32::FractionSize().0._State\ = \Posit32::FractionSize().0._State_6\) then 
                            \Posit32::FractionSize().0._State\ := \Posit32::FractionSize().0._State_5\;
                        end if;
                        
                    when \Posit32::FractionSize().0._State_7\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::FractionSize().0.conditionalf2eba7c459dd057c9270f346c2a9013399b4309fc21683746ef1be47061f03f1\ := to_unsigned(0, 32);
                        
                        if (\Posit32::FractionSize().0._State\ = \Posit32::FractionSize().0._State_7\) then 
                            \Posit32::FractionSize().0._State\ := \Posit32::FractionSize().0._State_5\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::FractionWithHiddenBit().0._StateMachine\: process (\Clock\) 
        Variable \Posit32::FractionWithHiddenBit().0._State\: \Posit32::FractionWithHiddenBit().0._States\ := \Posit32::FractionWithHiddenBit().0._State_0\;
        Variable \Posit32::FractionWithHiddenBit().0.this\: \Lombiq.Arithmetics.Posit32\;
        Variable \Posit32::FractionWithHiddenBit().0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::FractionWithHiddenBit().0.return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::FractionWithHiddenBit().0.num2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::FractionWithHiddenBit().0.conditionalec88d618fdb8d955a353066f43af5ab5cc70c1913e02ecac14c3590c5ee9802e\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::FractionWithHiddenBit().0.bits\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::FractionWithHiddenBit().0.binaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::FractionWithHiddenBit().0.binaryOperationResult.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::FractionWithHiddenBit().0.binaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::FractionWithHiddenBit().0.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::FractionWithHiddenBit().0.conditional7e2c70f465bbd6af6328e84460df8cc63262cd5e429e5f14f0c6d6c3620c3cea\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::FractionWithHiddenBit().0.binaryOperationResult.4\: boolean := false;
        Variable \Posit32::FractionWithHiddenBit().0.return.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::FractionWithHiddenBit().0._Finished\ <= false;
                \Posit32::FractionWithHiddenBit().0.return\ <= to_unsigned(0, 32);
                \Posit32::FractionWithHiddenBit().0.Posit32::FractionSize()._Started.0\ <= false;
                \Posit32::FractionWithHiddenBit().0.Posit32::SetOne(UInt32,UInt16).bits.parameter.Out.0\ <= to_unsigned(0, 32);
                \Posit32::FractionWithHiddenBit().0.Posit32::SetOne(UInt32,UInt16).index.parameter.Out.0\ <= to_unsigned(0, 16);
                \Posit32::FractionWithHiddenBit().0.Posit32::SetOne(UInt32,UInt16)._Started.0\ <= false;
                \Posit32::FractionWithHiddenBit().0._State\ := \Posit32::FractionWithHiddenBit().0._State_0\;
                \Posit32::FractionWithHiddenBit().0.num\ := to_unsigned(0, 32);
                \Posit32::FractionWithHiddenBit().0.return.0\ := to_unsigned(0, 32);
                \Posit32::FractionWithHiddenBit().0.num2\ := to_unsigned(0, 32);
                \Posit32::FractionWithHiddenBit().0.conditionalec88d618fdb8d955a353066f43af5ab5cc70c1913e02ecac14c3590c5ee9802e\ := to_unsigned(0, 32);
                \Posit32::FractionWithHiddenBit().0.bits\ := to_unsigned(0, 32);
                \Posit32::FractionWithHiddenBit().0.binaryOperationResult.0\ := to_signed(0, 32);
                \Posit32::FractionWithHiddenBit().0.binaryOperationResult.1\ := to_unsigned(0, 32);
                \Posit32::FractionWithHiddenBit().0.binaryOperationResult.2\ := to_signed(0, 32);
                \Posit32::FractionWithHiddenBit().0.binaryOperationResult.3\ := to_unsigned(0, 32);
                \Posit32::FractionWithHiddenBit().0.conditional7e2c70f465bbd6af6328e84460df8cc63262cd5e429e5f14f0c6d6c3620c3cea\ := to_unsigned(0, 32);
                \Posit32::FractionWithHiddenBit().0.binaryOperationResult.4\ := false;
                \Posit32::FractionWithHiddenBit().0.return.1\ := to_unsigned(0, 32);
            else 
                case \Posit32::FractionWithHiddenBit().0._State\ is 
                    when \Posit32::FractionWithHiddenBit().0._State_0\ => 
                        
                        
                        if (\Posit32::FractionWithHiddenBit().0._Started\ = true) then 
                            \Posit32::FractionWithHiddenBit().0._State\ := \Posit32::FractionWithHiddenBit().0._State_2\;
                        end if;
                        
                    when \Posit32::FractionWithHiddenBit().0._State_1\ => 
                        
                        
                        if (\Posit32::FractionWithHiddenBit().0._Started\ = true) then 
                            \Posit32::FractionWithHiddenBit().0._Finished\ <= true;
                        else 
                            \Posit32::FractionWithHiddenBit().0._Finished\ <= false;
                            \Posit32::FractionWithHiddenBit().0._State\ := \Posit32::FractionWithHiddenBit().0._State_0\;
                        end if;
                        
                    when \Posit32::FractionWithHiddenBit().0._State_2\ => 
                        \Posit32::FractionWithHiddenBit().0.this\ := \Posit32::FractionWithHiddenBit().0.this.parameter.In\;
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::FractionWithHiddenBit().0.Posit32::FractionSize().this.parameter.Out.0\ <= \Posit32::FractionWithHiddenBit().0.this\;
                        \Posit32::FractionWithHiddenBit().0.Posit32::FractionSize()._Started.0\ <= true;
                        \Posit32::FractionWithHiddenBit().0._State\ := \Posit32::FractionWithHiddenBit().0._State_3\;
                        
                    when \Posit32::FractionWithHiddenBit().0._State_3\ => 
                        
                        if (\Posit32::FractionWithHiddenBit().0.Posit32::FractionSize()._Started.0\ = \Posit32::FractionWithHiddenBit().0.Posit32::FractionSize()._Finished.0\) then 
                            \Posit32::FractionWithHiddenBit().0.Posit32::FractionSize()._Started.0\ <= false;
                            \Posit32::FractionWithHiddenBit().0.return.0\ := \Posit32::FractionWithHiddenBit().0.Posit32::FractionSize().return.0\;
                            \Posit32::FractionWithHiddenBit().0.num\ := \Posit32::FractionWithHiddenBit().0.return.0\;
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32::FractionWithHiddenBit().0.conditionalec88d618fdb8d955a353066f43af5ab5cc70c1913e02ecac14c3590c5ee9802e\ := to_unsigned(0, 32);
                            
                            
                            
                            \Posit32::FractionWithHiddenBit().0.num2\ := to_unsigned(0, 32);
                            
                            
                            
                            
                            
                            
                            \Posit32::FractionWithHiddenBit().0.binaryOperationResult.0\ := SmartResize(to_signed(32, 64) - signed(SmartResize((\Posit32::FractionWithHiddenBit().0.num\), 64)), 32);
                            \Posit32::FractionWithHiddenBit().0.binaryOperationResult.1\ := shift_left(to_unsigned(0, 32), to_integer(unsigned(SmartResize((\Posit32::FractionWithHiddenBit().0.binaryOperationResult.0\), 5))));
                            \Posit32::FractionWithHiddenBit().0._State\ := \Posit32::FractionWithHiddenBit().0._State_4\;
                        end if;
                        
                    when \Posit32::FractionWithHiddenBit().0._State_4\ => 
                        
                        \Posit32::FractionWithHiddenBit().0.binaryOperationResult.2\ := SmartResize(to_signed(32, 64) - signed(SmartResize((\Posit32::FractionWithHiddenBit().0.num\), 64)), 32);
                        \Posit32::FractionWithHiddenBit().0._State\ := \Posit32::FractionWithHiddenBit().0._State_5\;
                        
                    when \Posit32::FractionWithHiddenBit().0._State_5\ => 
                        
                        \Posit32::FractionWithHiddenBit().0.binaryOperationResult.3\ := shift_right(\Posit32::FractionWithHiddenBit().0.binaryOperationResult.1\, to_integer(unsigned(SmartResize((\Posit32::FractionWithHiddenBit().0.binaryOperationResult.2\), 5) and "11111")));
                        \Posit32::FractionWithHiddenBit().0.bits\ := \Posit32::FractionWithHiddenBit().0.binaryOperationResult.3\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::FractionWithHiddenBit().0._State\ := \Posit32::FractionWithHiddenBit().0._State_6\;
                        
                    when \Posit32::FractionWithHiddenBit().0._State_6\ => 
                        
                        \Posit32::FractionWithHiddenBit().0.binaryOperationResult.4\ := signed(SmartResize((\Posit32::FractionWithHiddenBit().0.num\), 64)) = to_signed(0, 64);

                        
                        
                        
                        

                        if ((\Posit32::FractionWithHiddenBit().0.binaryOperationResult.4\)) then 
                            \Posit32::FractionWithHiddenBit().0._State\ := \Posit32::FractionWithHiddenBit().0._State_8\;
                        else 
                            \Posit32::FractionWithHiddenBit().0._State\ := \Posit32::FractionWithHiddenBit().0._State_9\;
                        end if;
                        
                    when \Posit32::FractionWithHiddenBit().0._State_7\ => 
                        
                        
                        
                        
                        \Posit32::FractionWithHiddenBit().0.return\ <= \Posit32::FractionWithHiddenBit().0.conditional7e2c70f465bbd6af6328e84460df8cc63262cd5e429e5f14f0c6d6c3620c3cea\;
                        \Posit32::FractionWithHiddenBit().0._State\ := \Posit32::FractionWithHiddenBit().0._State_1\;
                        
                    when \Posit32::FractionWithHiddenBit().0._State_8\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::FractionWithHiddenBit().0.conditional7e2c70f465bbd6af6328e84460df8cc63262cd5e429e5f14f0c6d6c3620c3cea\ := to_unsigned(1, 32);
                        
                        if (\Posit32::FractionWithHiddenBit().0._State\ = \Posit32::FractionWithHiddenBit().0._State_8\) then 
                            \Posit32::FractionWithHiddenBit().0._State\ := \Posit32::FractionWithHiddenBit().0._State_7\;
                        end if;
                        
                    when \Posit32::FractionWithHiddenBit().0._State_9\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::FractionWithHiddenBit().0.Posit32::SetOne(UInt32,UInt16).this.parameter.Out.0\ <= \Posit32::FractionWithHiddenBit().0.this\;
                        \Posit32::FractionWithHiddenBit().0.Posit32::SetOne(UInt32,UInt16).bits.parameter.Out.0\ <= \Posit32::FractionWithHiddenBit().0.bits\;
                        \Posit32::FractionWithHiddenBit().0.Posit32::SetOne(UInt32,UInt16).index.parameter.Out.0\ <= SmartResize(\Posit32::FractionWithHiddenBit().0.num\, 16);
                        \Posit32::FractionWithHiddenBit().0.Posit32::SetOne(UInt32,UInt16)._Started.0\ <= true;
                        \Posit32::FractionWithHiddenBit().0._State\ := \Posit32::FractionWithHiddenBit().0._State_10\;
                        
                    when \Posit32::FractionWithHiddenBit().0._State_10\ => 
                        
                        if (\Posit32::FractionWithHiddenBit().0.Posit32::SetOne(UInt32,UInt16)._Started.0\ = \Posit32::FractionWithHiddenBit().0.Posit32::SetOne(UInt32,UInt16)._Finished.0\) then 
                            \Posit32::FractionWithHiddenBit().0.Posit32::SetOne(UInt32,UInt16)._Started.0\ <= false;
                            \Posit32::FractionWithHiddenBit().0.return.1\ := \Posit32::FractionWithHiddenBit().0.Posit32::SetOne(UInt32,UInt16).return.0\;
                            \Posit32::FractionWithHiddenBit().0.conditional7e2c70f465bbd6af6328e84460df8cc63262cd5e429e5f14f0c6d6c3620c3cea\ := \Posit32::FractionWithHiddenBit().0.return.1\;
                            
                            if (\Posit32::FractionWithHiddenBit().0._State\ = \Posit32::FractionWithHiddenBit().0._State_10\) then 
                                \Posit32::FractionWithHiddenBit().0._State\ := \Posit32::FractionWithHiddenBit().0._State_7\;
                            end if;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::GetMostSignificantOnePosition(UInt32).0._StateMachine\: process (\Clock\) 
        Variable \Posit32::GetMostSignificantOnePosition(UInt32).0._State\: \Posit32::GetMostSignificantOnePosition(UInt32).0._States\ := \Posit32::GetMostSignificantOnePosition(UInt32).0._State_0\;
        Variable \Posit32::GetMostSignificantOnePosition(UInt32).0.bits\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::GetMostSignificantOnePosition(UInt32).0.b\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::GetMostSignificantOnePosition(UInt32).0.binaryOperationResult.0\: boolean := false;
        Variable \Posit32::GetMostSignificantOnePosition(UInt32).0.binaryOperationResult.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::GetMostSignificantOnePosition(UInt32).0.binaryOperationResult.2\: unsigned(7 downto 0) := to_unsigned(0, 8);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::GetMostSignificantOnePosition(UInt32).0._Finished\ <= false;
                \Posit32::GetMostSignificantOnePosition(UInt32).0.return\ <= to_unsigned(0, 8);
                \Posit32::GetMostSignificantOnePosition(UInt32).0._State\ := \Posit32::GetMostSignificantOnePosition(UInt32).0._State_0\;
                \Posit32::GetMostSignificantOnePosition(UInt32).0.bits\ := to_unsigned(0, 32);
                \Posit32::GetMostSignificantOnePosition(UInt32).0.b\ := to_unsigned(0, 8);
                \Posit32::GetMostSignificantOnePosition(UInt32).0.binaryOperationResult.0\ := false;
                \Posit32::GetMostSignificantOnePosition(UInt32).0.binaryOperationResult.1\ := to_unsigned(0, 32);
                \Posit32::GetMostSignificantOnePosition(UInt32).0.binaryOperationResult.2\ := to_unsigned(0, 8);
            else 
                case \Posit32::GetMostSignificantOnePosition(UInt32).0._State\ is 
                    when \Posit32::GetMostSignificantOnePosition(UInt32).0._State_0\ => 
                        
                        
                        if (\Posit32::GetMostSignificantOnePosition(UInt32).0._Started\ = true) then 
                            \Posit32::GetMostSignificantOnePosition(UInt32).0._State\ := \Posit32::GetMostSignificantOnePosition(UInt32).0._State_2\;
                        end if;
                        
                    when \Posit32::GetMostSignificantOnePosition(UInt32).0._State_1\ => 
                        
                        
                        if (\Posit32::GetMostSignificantOnePosition(UInt32).0._Started\ = true) then 
                            \Posit32::GetMostSignificantOnePosition(UInt32).0._Finished\ <= true;
                        else 
                            \Posit32::GetMostSignificantOnePosition(UInt32).0._Finished\ <= false;
                            \Posit32::GetMostSignificantOnePosition(UInt32).0._State\ := \Posit32::GetMostSignificantOnePosition(UInt32).0._State_0\;
                        end if;
                        
                    when \Posit32::GetMostSignificantOnePosition(UInt32).0._State_2\ => 
                        \Posit32::GetMostSignificantOnePosition(UInt32).0.bits\ := \Posit32::GetMostSignificantOnePosition(UInt32).0.bits.parameter.In\;
                        
                        
                        
                        
                        
                        
                        \Posit32::GetMostSignificantOnePosition(UInt32).0.b\ := SmartResize(unsigned(to_signed(0, 32)), 8);
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::GetMostSignificantOnePosition(UInt32).0._State\ := \Posit32::GetMostSignificantOnePosition(UInt32).0._State_3\;
                        
                    when \Posit32::GetMostSignificantOnePosition(UInt32).0._State_3\ => 
                        
                        
                        \Posit32::GetMostSignificantOnePosition(UInt32).0.binaryOperationResult.0\ := signed(SmartResize((\Posit32::GetMostSignificantOnePosition(UInt32).0.bits\), 64)) /= to_signed(0, 64);
                        if (\Posit32::GetMostSignificantOnePosition(UInt32).0.binaryOperationResult.0\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32::GetMostSignificantOnePosition(UInt32).0.binaryOperationResult.1\ := shift_right(\Posit32::GetMostSignificantOnePosition(UInt32).0.bits\, to_integer(unsigned(SmartResize(to_signed(1, 32), 5) and "11111")));
                            \Posit32::GetMostSignificantOnePosition(UInt32).0.bits\ := \Posit32::GetMostSignificantOnePosition(UInt32).0.binaryOperationResult.1\;
                            
                            
                            
                            \Posit32::GetMostSignificantOnePosition(UInt32).0._State\ := \Posit32::GetMostSignificantOnePosition(UInt32).0._State_5\;
                        else 
                            \Posit32::GetMostSignificantOnePosition(UInt32).0._State\ := \Posit32::GetMostSignificantOnePosition(UInt32).0._State_4\;
                        end if;
                        
                    when \Posit32::GetMostSignificantOnePosition(UInt32).0._State_4\ => 
                        
                        
                        
                        
                        \Posit32::GetMostSignificantOnePosition(UInt32).0.return\ <= \Posit32::GetMostSignificantOnePosition(UInt32).0.b\;
                        \Posit32::GetMostSignificantOnePosition(UInt32).0._State\ := \Posit32::GetMostSignificantOnePosition(UInt32).0._State_1\;
                        
                    when \Posit32::GetMostSignificantOnePosition(UInt32).0._State_5\ => 
                        
                        \Posit32::GetMostSignificantOnePosition(UInt32).0.binaryOperationResult.2\ := SmartResize(unsigned(signed(SmartResize((\Posit32::GetMostSignificantOnePosition(UInt32).0.b\), 32)) + to_signed(1, 32)), 8);
                        \Posit32::GetMostSignificantOnePosition(UInt32).0.b\ := (\Posit32::GetMostSignificantOnePosition(UInt32).0.binaryOperationResult.2\);
                        
                        if (\Posit32::GetMostSignificantOnePosition(UInt32).0._State\ = \Posit32::GetMostSignificantOnePosition(UInt32).0._State_5\) then 
                            \Posit32::GetMostSignificantOnePosition(UInt32).0._State\ := \Posit32::GetMostSignificantOnePosition(UInt32).0._State_3\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::SetOne(UInt32,UInt16).0._StateMachine\: process (\Clock\) 
        Variable \Posit32::SetOne(UInt32,UInt16).0._State\: \Posit32::SetOne(UInt32,UInt16).0._States\ := \Posit32::SetOne(UInt32,UInt16).0._State_0\;
        Variable \Posit32::SetOne(UInt32,UInt16).0.this\: \Lombiq.Arithmetics.Posit32\;
        Variable \Posit32::SetOne(UInt32,UInt16).0.bits\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::SetOne(UInt32,UInt16).0.index\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Posit32::SetOne(UInt32,UInt16).0.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::SetOne(UInt32,UInt16).0.binaryOperationResult.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::SetOne(UInt32,UInt16).0._Finished\ <= false;
                \Posit32::SetOne(UInt32,UInt16).0.return\ <= to_unsigned(0, 32);
                \Posit32::SetOne(UInt32,UInt16).0._State\ := \Posit32::SetOne(UInt32,UInt16).0._State_0\;
                \Posit32::SetOne(UInt32,UInt16).0.bits\ := to_unsigned(0, 32);
                \Posit32::SetOne(UInt32,UInt16).0.index\ := to_unsigned(0, 16);
                \Posit32::SetOne(UInt32,UInt16).0.binaryOperationResult.0\ := to_unsigned(0, 32);
                \Posit32::SetOne(UInt32,UInt16).0.binaryOperationResult.1\ := to_unsigned(0, 32);
            else 
                case \Posit32::SetOne(UInt32,UInt16).0._State\ is 
                    when \Posit32::SetOne(UInt32,UInt16).0._State_0\ => 
                        
                        
                        if (\Posit32::SetOne(UInt32,UInt16).0._Started\ = true) then 
                            \Posit32::SetOne(UInt32,UInt16).0._State\ := \Posit32::SetOne(UInt32,UInt16).0._State_2\;
                        end if;
                        
                    when \Posit32::SetOne(UInt32,UInt16).0._State_1\ => 
                        
                        
                        if (\Posit32::SetOne(UInt32,UInt16).0._Started\ = true) then 
                            \Posit32::SetOne(UInt32,UInt16).0._Finished\ <= true;
                        else 
                            \Posit32::SetOne(UInt32,UInt16).0._Finished\ <= false;
                            \Posit32::SetOne(UInt32,UInt16).0._State\ := \Posit32::SetOne(UInt32,UInt16).0._State_0\;
                        end if;
                        
                    when \Posit32::SetOne(UInt32,UInt16).0._State_2\ => 
                        \Posit32::SetOne(UInt32,UInt16).0.this\ := \Posit32::SetOne(UInt32,UInt16).0.this.parameter.In\;
                        \Posit32::SetOne(UInt32,UInt16).0.bits\ := \Posit32::SetOne(UInt32,UInt16).0.bits.parameter.In\;
                        \Posit32::SetOne(UInt32,UInt16).0.index\ := \Posit32::SetOne(UInt32,UInt16).0.index.parameter.In\;
                        
                        
                        
                        \Posit32::SetOne(UInt32,UInt16).0.binaryOperationResult.0\ := unsigned(shift_left(to_signed(1, 32), to_integer(unsigned(SmartResize(signed(SmartResize(\Posit32::SetOne(UInt32,UInt16).0.index\, 32)), 5)))));
                        \Posit32::SetOne(UInt32,UInt16).0.binaryOperationResult.1\ := \Posit32::SetOne(UInt32,UInt16).0.bits\ or (\Posit32::SetOne(UInt32,UInt16).0.binaryOperationResult.0\);
                        \Posit32::SetOne(UInt32,UInt16).0.return\ <= \Posit32::SetOne(UInt32,UInt16).0.binaryOperationResult.1\;
                        \Posit32::SetOne(UInt32,UInt16).0._State\ := \Posit32::SetOne(UInt32,UInt16).0._State_1\;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::SetZero(UInt32,UInt16).0._StateMachine\: process (\Clock\) 
        Variable \Posit32::SetZero(UInt32,UInt16).0._State\: \Posit32::SetZero(UInt32,UInt16).0._States\ := \Posit32::SetZero(UInt32,UInt16).0._State_0\;
        Variable \Posit32::SetZero(UInt32,UInt16).0.bits\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::SetZero(UInt32,UInt16).0.index\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Posit32::SetZero(UInt32,UInt16).0.binaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::SetZero(UInt32,UInt16).0.unaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::SetZero(UInt32,UInt16).0.binaryOperationResult.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::SetZero(UInt32,UInt16).0._Finished\ <= false;
                \Posit32::SetZero(UInt32,UInt16).0.return\ <= to_unsigned(0, 32);
                \Posit32::SetZero(UInt32,UInt16).0._State\ := \Posit32::SetZero(UInt32,UInt16).0._State_0\;
                \Posit32::SetZero(UInt32,UInt16).0.bits\ := to_unsigned(0, 32);
                \Posit32::SetZero(UInt32,UInt16).0.index\ := to_unsigned(0, 16);
                \Posit32::SetZero(UInt32,UInt16).0.binaryOperationResult.0\ := to_signed(0, 32);
                \Posit32::SetZero(UInt32,UInt16).0.unaryOperationResult.0\ := to_signed(0, 32);
                \Posit32::SetZero(UInt32,UInt16).0.binaryOperationResult.1\ := to_unsigned(0, 32);
            else 
                case \Posit32::SetZero(UInt32,UInt16).0._State\ is 
                    when \Posit32::SetZero(UInt32,UInt16).0._State_0\ => 
                        
                        
                        if (\Posit32::SetZero(UInt32,UInt16).0._Started\ = true) then 
                            \Posit32::SetZero(UInt32,UInt16).0._State\ := \Posit32::SetZero(UInt32,UInt16).0._State_2\;
                        end if;
                        
                    when \Posit32::SetZero(UInt32,UInt16).0._State_1\ => 
                        
                        
                        if (\Posit32::SetZero(UInt32,UInt16).0._Started\ = true) then 
                            \Posit32::SetZero(UInt32,UInt16).0._Finished\ <= true;
                        else 
                            \Posit32::SetZero(UInt32,UInt16).0._Finished\ <= false;
                            \Posit32::SetZero(UInt32,UInt16).0._State\ := \Posit32::SetZero(UInt32,UInt16).0._State_0\;
                        end if;
                        
                    when \Posit32::SetZero(UInt32,UInt16).0._State_2\ => 
                        \Posit32::SetZero(UInt32,UInt16).0.bits\ := \Posit32::SetZero(UInt32,UInt16).0.bits.parameter.In\;
                        \Posit32::SetZero(UInt32,UInt16).0.index\ := \Posit32::SetZero(UInt32,UInt16).0.index.parameter.In\;
                        
                        
                        
                        \Posit32::SetZero(UInt32,UInt16).0.binaryOperationResult.0\ := shift_left(to_signed(1, 32), to_integer(unsigned(SmartResize(signed(SmartResize(\Posit32::SetZero(UInt32,UInt16).0.index\, 32)), 5))));
                        \Posit32::SetZero(UInt32,UInt16).0.unaryOperationResult.0\ := not((\Posit32::SetZero(UInt32,UInt16).0.binaryOperationResult.0\));
                        \Posit32::SetZero(UInt32,UInt16).0.binaryOperationResult.1\ := \Posit32::SetZero(UInt32,UInt16).0.bits\ and unsigned((\Posit32::SetZero(UInt32,UInt16).0.unaryOperationResult.0\));
                        \Posit32::SetZero(UInt32,UInt16).0.return\ <= \Posit32::SetZero(UInt32,UInt16).0.binaryOperationResult.1\;
                        \Posit32::SetZero(UInt32,UInt16).0._State\ := \Posit32::SetZero(UInt32,UInt16).0._State_1\;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::LengthOfRunOfBits(UInt32,Byte).0._StateMachine\: process (\Clock\) 
        Variable \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State\: \Posit32::LengthOfRunOfBits(UInt32,Byte).0._States\ := \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_0\;
        Variable \Posit32::LengthOfRunOfBits(UInt32,Byte).0.bits\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::LengthOfRunOfBits(UInt32,Byte).0.startingPosition\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::LengthOfRunOfBits(UInt32,Byte).0.b\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::LengthOfRunOfBits(UInt32,Byte).0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::LengthOfRunOfBits(UInt32,Byte).0.num2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.4\: boolean := false;
        Variable \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.5\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.6\: boolean := false;
        Variable \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.7\: boolean := false;
        Variable \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.8\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.9\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.10\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::LengthOfRunOfBits(UInt32,Byte).0._Finished\ <= false;
                \Posit32::LengthOfRunOfBits(UInt32,Byte).0.return\ <= to_unsigned(0, 8);
                \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State\ := \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_0\;
                \Posit32::LengthOfRunOfBits(UInt32,Byte).0.bits\ := to_unsigned(0, 32);
                \Posit32::LengthOfRunOfBits(UInt32,Byte).0.startingPosition\ := to_unsigned(0, 8);
                \Posit32::LengthOfRunOfBits(UInt32,Byte).0.b\ := to_unsigned(0, 8);
                \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.0\ := to_unsigned(0, 32);
                \Posit32::LengthOfRunOfBits(UInt32,Byte).0.num\ := to_unsigned(0, 32);
                \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.1\ := to_unsigned(0, 32);
                \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.2\ := to_unsigned(0, 32);
                \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.3\ := to_unsigned(0, 32);
                \Posit32::LengthOfRunOfBits(UInt32,Byte).0.num2\ := to_signed(0, 32);
                \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.4\ := false;
                \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.5\ := to_unsigned(0, 32);
                \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.6\ := false;
                \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.7\ := false;
                \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.8\ := to_unsigned(0, 32);
                \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.9\ := to_unsigned(0, 8);
                \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.10\ := to_signed(0, 32);
            else 
                case \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State\ is 
                    when \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_0\ => 
                        
                        
                        if (\Posit32::LengthOfRunOfBits(UInt32,Byte).0._Started\ = true) then 
                            \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State\ := \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_2\;
                        end if;
                        
                    when \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_1\ => 
                        
                        
                        if (\Posit32::LengthOfRunOfBits(UInt32,Byte).0._Started\ = true) then 
                            \Posit32::LengthOfRunOfBits(UInt32,Byte).0._Finished\ <= true;
                        else 
                            \Posit32::LengthOfRunOfBits(UInt32,Byte).0._Finished\ <= false;
                            \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State\ := \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_0\;
                        end if;
                        
                    when \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_2\ => 
                        \Posit32::LengthOfRunOfBits(UInt32,Byte).0.bits\ := \Posit32::LengthOfRunOfBits(UInt32,Byte).0.bits.parameter.In\;
                        \Posit32::LengthOfRunOfBits(UInt32,Byte).0.startingPosition\ := \Posit32::LengthOfRunOfBits(UInt32,Byte).0.startingPosition.parameter.In\;
                        
                        
                        
                        
                        
                        
                        \Posit32::LengthOfRunOfBits(UInt32,Byte).0.b\ := SmartResize(unsigned(to_signed(1, 32)), 8);
                        
                        
                        
                        \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.0\ := shift_left(\Posit32::LengthOfRunOfBits(UInt32,Byte).0.bits\, to_integer(unsigned(SmartResize(to_signed(1, 32), 5))));
                        \Posit32::LengthOfRunOfBits(UInt32,Byte).0.bits\ := \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.0\;
                        
                        
                        
                        
                        
                        
                        \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.1\ := shift_right(\Posit32::LengthOfRunOfBits(UInt32,Byte).0.bits\, to_integer(unsigned(SmartResize(to_signed(31, 32), 5) and "11111")));
                        \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.2\ := (\Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.1\) and to_unsigned(1, 32);
                        \Posit32::LengthOfRunOfBits(UInt32,Byte).0.num\ := \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.2\;
                        
                        
                        
                        \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.3\ := shift_left(\Posit32::LengthOfRunOfBits(UInt32,Byte).0.bits\, to_integer(unsigned(SmartResize(to_signed(1, 32), 5))));
                        \Posit32::LengthOfRunOfBits(UInt32,Byte).0.bits\ := \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.3\;
                        
                        
                        
                        
                        
                        
                        \Posit32::LengthOfRunOfBits(UInt32,Byte).0.num2\ := to_signed(0, 32);
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State\ := \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_3\;
                        
                    when \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_3\ => 
                        
                        
                        \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.4\ := (\Posit32::LengthOfRunOfBits(UInt32,Byte).0.num2\) < signed(SmartResize((\Posit32::LengthOfRunOfBits(UInt32,Byte).0.startingPosition\), 32));
                        \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.5\ := shift_right(\Posit32::LengthOfRunOfBits(UInt32,Byte).0.bits\, to_integer(unsigned(SmartResize(to_signed(31, 32), 5) and "11111")));
                        \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State\ := \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_5\;
                        
                    when \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_4\ => 
                        
                        
                        
                        
                        \Posit32::LengthOfRunOfBits(UInt32,Byte).0.return\ <= \Posit32::LengthOfRunOfBits(UInt32,Byte).0.b\;
                        \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State\ := \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_1\;
                        
                    when \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_5\ => 
                        
                        \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.6\ := \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.5\ = \Posit32::LengthOfRunOfBits(UInt32,Byte).0.num\;
                        \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.7\ := \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.4\ and \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.6\;
                        if (\Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.7\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.8\ := shift_left(\Posit32::LengthOfRunOfBits(UInt32,Byte).0.bits\, to_integer(unsigned(SmartResize(to_signed(1, 32), 5))));
                            \Posit32::LengthOfRunOfBits(UInt32,Byte).0.bits\ := \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.8\;
                            
                            
                            
                            \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State\ := \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_6\;
                        else 
                            \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State\ := \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_4\;
                        end if;
                        
                    when \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_6\ => 
                        
                        \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.9\ := SmartResize(unsigned(signed(SmartResize((\Posit32::LengthOfRunOfBits(UInt32,Byte).0.b\), 32)) + to_signed(1, 32)), 8);
                        \Posit32::LengthOfRunOfBits(UInt32,Byte).0.b\ := (\Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.9\);
                        
                        
                        
                        \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.10\ := \Posit32::LengthOfRunOfBits(UInt32,Byte).0.num2\ + to_signed(1, 32);
                        \Posit32::LengthOfRunOfBits(UInt32,Byte).0.num2\ := \Posit32::LengthOfRunOfBits(UInt32,Byte).0.binaryOperationResult.10\;
                        
                        if (\Posit32::LengthOfRunOfBits(UInt32,Byte).0._State\ = \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_6\) then 
                            \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State\ := \Posit32::LengthOfRunOfBits(UInt32,Byte).0._State_3\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::GetTwosComplement(UInt32).0._StateMachine\: process (\Clock\) 
        Variable \Posit32::GetTwosComplement(UInt32).0._State\: \Posit32::GetTwosComplement(UInt32).0._States\ := \Posit32::GetTwosComplement(UInt32).0._State_0\;
        Variable \Posit32::GetTwosComplement(UInt32).0.bits\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::GetTwosComplement(UInt32).0.unaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::GetTwosComplement(UInt32).0.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::GetTwosComplement(UInt32).0._Finished\ <= false;
                \Posit32::GetTwosComplement(UInt32).0.return\ <= to_unsigned(0, 32);
                \Posit32::GetTwosComplement(UInt32).0._State\ := \Posit32::GetTwosComplement(UInt32).0._State_0\;
                \Posit32::GetTwosComplement(UInt32).0.bits\ := to_unsigned(0, 32);
                \Posit32::GetTwosComplement(UInt32).0.unaryOperationResult.0\ := to_unsigned(0, 32);
                \Posit32::GetTwosComplement(UInt32).0.binaryOperationResult.0\ := to_unsigned(0, 32);
            else 
                case \Posit32::GetTwosComplement(UInt32).0._State\ is 
                    when \Posit32::GetTwosComplement(UInt32).0._State_0\ => 
                        
                        
                        if (\Posit32::GetTwosComplement(UInt32).0._Started\ = true) then 
                            \Posit32::GetTwosComplement(UInt32).0._State\ := \Posit32::GetTwosComplement(UInt32).0._State_2\;
                        end if;
                        
                    when \Posit32::GetTwosComplement(UInt32).0._State_1\ => 
                        
                        
                        if (\Posit32::GetTwosComplement(UInt32).0._Started\ = true) then 
                            \Posit32::GetTwosComplement(UInt32).0._Finished\ <= true;
                        else 
                            \Posit32::GetTwosComplement(UInt32).0._Finished\ <= false;
                            \Posit32::GetTwosComplement(UInt32).0._State\ := \Posit32::GetTwosComplement(UInt32).0._State_0\;
                        end if;
                        
                    when \Posit32::GetTwosComplement(UInt32).0._State_2\ => 
                        \Posit32::GetTwosComplement(UInt32).0.bits\ := \Posit32::GetTwosComplement(UInt32).0.bits.parameter.In\;
                        
                        
                        
                        \Posit32::GetTwosComplement(UInt32).0.unaryOperationResult.0\ := not(\Posit32::GetTwosComplement(UInt32).0.bits\);
                        \Posit32::GetTwosComplement(UInt32).0.binaryOperationResult.0\ := SmartResize(unsigned(signed(SmartResize((\Posit32::GetTwosComplement(UInt32).0.unaryOperationResult.0\), 64)) + to_signed(1, 64)), 32);
                        \Posit32::GetTwosComplement(UInt32).0.return\ <= (\Posit32::GetTwosComplement(UInt32).0.binaryOperationResult.0\);
                        \Posit32::GetTwosComplement(UInt32).0._State\ := \Posit32::GetTwosComplement(UInt32).0._State_1\;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::FusedSum(Posit32[],Quire).0._StateMachine\: process (\Clock\) 
        Variable \Posit32::FusedSum(Posit32[],Quire).0._State\: \Posit32::FusedSum(Posit32[],Quire).0._States\ := \Posit32::FusedSum(Posit32[],Quire).0._State_0\;
        Variable \Posit32::FusedSum(Posit32[],Quire).0.posits\: \Lombiq.Arithmetics.Posit32_Array\(0 to 159);
        Variable \Posit32::FusedSum(Posit32[],Quire).0.startingValue\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::FusedSum(Posit32[],Quire).0.quire\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::FusedSum(Posit32[],Quire).0.objectcca0dec009ae8ed2326a07122a465f3ec1a2db6344ea5f25f4320f84fc89c011\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::FusedSum(Posit32[],Quire).0.return.0\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::FusedSum(Posit32[],Quire).0.return.1\: boolean := false;
        Variable \Posit32::FusedSum(Posit32[],Quire).0.num\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::FusedSum(Posit32[],Quire).0.binaryOperationResult.0\: boolean := false;
        Variable \Posit32::FusedSum(Posit32[],Quire).0.return.2\: boolean := false;
        Variable \Posit32::FusedSum(Posit32[],Quire).0.return.3\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::FusedSum(Posit32[],Quire).0.return.4\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::FusedSum(Posit32[],Quire).0.binaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::FusedSum(Posit32[],Quire).0._Finished\ <= false;
                \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).firstSegment.parameter.Out.0\ <= to_unsigned(0, 32);
                \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Started.0\ <= false;
                \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\ <= to_signed(0, 32);
                \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ <= false;
                \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire)._Started.0\ <= false;
                \Posit32::FusedSum(Posit32[],Quire).0.Posit32::IsNaN()._Started.0\ <= false;
                \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Started.0\ <= false;
                \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\ <= false;
                \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_0\;
                \Posit32::FusedSum(Posit32[],Quire).0.return.1\ := false;
                \Posit32::FusedSum(Posit32[],Quire).0.num\ := to_signed(0, 32);
                \Posit32::FusedSum(Posit32[],Quire).0.binaryOperationResult.0\ := false;
                \Posit32::FusedSum(Posit32[],Quire).0.return.2\ := false;
                \Posit32::FusedSum(Posit32[],Quire).0.binaryOperationResult.1\ := to_signed(0, 32);
            else 
                case \Posit32::FusedSum(Posit32[],Quire).0._State\ is 
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_0\ => 
                        
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0._Started\ = true) then 
                            \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_2\;
                        end if;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_1\ => 
                        
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0._Started\ = true) then 
                            \Posit32::FusedSum(Posit32[],Quire).0._Finished\ <= true;
                        else 
                            \Posit32::FusedSum(Posit32[],Quire).0._Finished\ <= false;
                            \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_0\;
                        end if;
                        
                        \Posit32::FusedSum(Posit32[],Quire).0.posits.parameter.Out\ <= \Posit32::FusedSum(Posit32[],Quire).0.posits\;
                        \Posit32::FusedSum(Posit32[],Quire).0.startingValue.parameter.Out\ <= \Posit32::FusedSum(Posit32[],Quire).0.startingValue\;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_2\ => 
                        \Posit32::FusedSum(Posit32[],Quire).0.posits\ := \Posit32::FusedSum(Posit32[],Quire).0.posits.parameter.In\;
                        \Posit32::FusedSum(Posit32[],Quire).0.startingValue\ := \Posit32::FusedSum(Posit32[],Quire).0.startingValue.parameter.In\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::FusedSum(Posit32[],Quire).0.objectcca0dec009ae8ed2326a07122a465f3ec1a2db6344ea5f25f4320f84fc89c011\.\IsNull\ := false;
                        \Posit32::FusedSum(Posit32[],Quire).0.objectcca0dec009ae8ed2326a07122a465f3ec1a2db6344ea5f25f4320f84fc89c011\.\Size\ := to_unsigned(0, 16);
                        \Posit32::FusedSum(Posit32[],Quire).0.objectcca0dec009ae8ed2326a07122a465f3ec1a2db6344ea5f25f4320f84fc89c011\.\SegmentCount\ := to_unsigned(0, 16);
                        \Posit32::FusedSum(Posit32[],Quire).0.objectcca0dec009ae8ed2326a07122a465f3ec1a2db6344ea5f25f4320f84fc89c011\.\Segments\ := (others => to_unsigned(0, 64));
                        
                        
                        \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).this.parameter.Out.0\ <= \Posit32::FusedSum(Posit32[],Quire).0.objectcca0dec009ae8ed2326a07122a465f3ec1a2db6344ea5f25f4320f84fc89c011\;
                        \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).firstSegment.parameter.Out.0\ <= to_unsigned(1, 32);
                        \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).size.parameter.Out.0\ <= SmartResize(unsigned(to_signed(512, 32)), 16);
                        \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Started.0\ <= true;
                        \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_3\;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_3\ => 
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Started.0\ = \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Finished.0\) then 
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Started.0\ <= false;
                            \Posit32::FusedSum(Posit32[],Quire).0.objectcca0dec009ae8ed2326a07122a465f3ec1a2db6344ea5f25f4320f84fc89c011\ := \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).this.parameter.In.0\;
                            
                            
                            
                            
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.Out.0\ <= \Posit32::FusedSum(Posit32[],Quire).0.objectcca0dec009ae8ed2326a07122a465f3ec1a2db6344ea5f25f4320f84fc89c011\;
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\ <= to_signed(511, 32);
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ <= true;
                            \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_4\;
                        end if;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_4\ => 
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ = \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\) then 
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ <= false;
                            \Posit32::FusedSum(Posit32[],Quire).0.return.0\ := \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).return.0\;
                            \Posit32::FusedSum(Posit32[],Quire).0.objectcca0dec009ae8ed2326a07122a465f3ec1a2db6344ea5f25f4320f84fc89c011\ := \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.In.0\;
                            \Posit32::FusedSum(Posit32[],Quire).0.quire\ := \Posit32::FusedSum(Posit32[],Quire).0.return.0\;
                            
                            
                            
                            
                            
                            
                            \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).left.parameter.Out.0\ <= \Posit32::FusedSum(Posit32[],Quire).0.startingValue\;
                            \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).right.parameter.Out.0\ <= \Posit32::FusedSum(Posit32[],Quire).0.quire\;
                            \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire)._Started.0\ <= true;
                            \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_5\;
                        end if;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_5\ => 
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire)._Started.0\ = \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire)._Finished.0\) then 
                            \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire)._Started.0\ <= false;
                            \Posit32::FusedSum(Posit32[],Quire).0.return.1\ := \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).return.0\;
                            \Posit32::FusedSum(Posit32[],Quire).0.startingValue\ := \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).left.parameter.In.0\;
                            \Posit32::FusedSum(Posit32[],Quire).0.quire\ := \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).right.parameter.In.0\;

                            
                            
                            

                            if (\Posit32::FusedSum(Posit32[],Quire).0.return.1\) then 
                                \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_7\;
                            else 
                                
                                \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_6\;
                            end if;
                        end if;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_6\ => 
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::FusedSum(Posit32[],Quire).0.num\ := to_signed(0, 32);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_8\;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_7\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::FusedSum(Posit32[],Quire).0.return\ <= \Posit32::FusedSum(Posit32[],Quire).0.quire\;
                        \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_1\;
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0._State\ = \Posit32::FusedSum(Posit32[],Quire).0._State_7\) then 
                            \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_6\;
                        end if;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_8\ => 
                        
                        
                        \Posit32::FusedSum(Posit32[],Quire).0.binaryOperationResult.0\ := \Posit32::FusedSum(Posit32[],Quire).0.num\ < to_signed(160, 32);
                        if (\Posit32::FusedSum(Posit32[],Quire).0.binaryOperationResult.0\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32::FusedSum(Posit32[],Quire).0.Posit32::IsNaN().this.parameter.Out.0\ <= \Posit32::FusedSum(Posit32[],Quire).0.posits\(to_integer(\Posit32::FusedSum(Posit32[],Quire).0.num\));
                            \Posit32::FusedSum(Posit32[],Quire).0.Posit32::IsNaN()._Started.0\ <= true;
                            \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_10\;
                        else 
                            \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_9\;
                        end if;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_9\ => 
                        
                        
                        
                        
                        \Posit32::FusedSum(Posit32[],Quire).0.return\ <= \Posit32::FusedSum(Posit32[],Quire).0.startingValue\;
                        \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_1\;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_10\ => 
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Posit32::IsNaN()._Started.0\ = \Posit32::FusedSum(Posit32[],Quire).0.Posit32::IsNaN()._Finished.0\) then 
                            \Posit32::FusedSum(Posit32[],Quire).0.Posit32::IsNaN()._Started.0\ <= false;
                            \Posit32::FusedSum(Posit32[],Quire).0.return.2\ := \Posit32::FusedSum(Posit32[],Quire).0.Posit32::IsNaN().return.0\;

                            
                            
                            

                            if (\Posit32::FusedSum(Posit32[],Quire).0.return.2\) then 
                                \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_12\;
                            else 
                                
                                \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_11\;
                            end if;
                        end if;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_11\ => 
                        
                        
                        
                        
                        
                        \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32).x.parameter.Out.0\ <= \Posit32::FusedSum(Posit32[],Quire).0.posits\(to_integer(\Posit32::FusedSum(Posit32[],Quire).0.num\));
                        \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Started.0\ <= true;
                        \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_13\;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_12\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::FusedSum(Posit32[],Quire).0.return\ <= \Posit32::FusedSum(Posit32[],Quire).0.quire\;
                        \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_1\;
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0._State\ = \Posit32::FusedSum(Posit32[],Quire).0._State_12\) then 
                            \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_11\;
                        end if;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_13\ => 
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Started.0\ = \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\) then 
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Started.0\ <= false;
                            \Posit32::FusedSum(Posit32[],Quire).0.return.3\ := \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32).return.0\;
                            
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.Out.0\ <= \Posit32::FusedSum(Posit32[],Quire).0.startingValue\;
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.Out.0\ <= \Posit32::FusedSum(Posit32[],Quire).0.return.3\;
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\ <= true;
                            \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_14\;
                        end if;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_14\ => 
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\ = \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\) then 
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\ <= false;
                            \Posit32::FusedSum(Posit32[],Quire).0.return.4\ := \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).return.0\;
                            \Posit32::FusedSum(Posit32[],Quire).0.startingValue\ := \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.In.0\;
                            \Posit32::FusedSum(Posit32[],Quire).0.return.3\ := \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.In.0\;
                            \Posit32::FusedSum(Posit32[],Quire).0.startingValue\ := \Posit32::FusedSum(Posit32[],Quire).0.return.4\;
                            
                            
                            
                            \Posit32::FusedSum(Posit32[],Quire).0.binaryOperationResult.1\ := \Posit32::FusedSum(Posit32[],Quire).0.num\ + to_signed(1, 32);
                            \Posit32::FusedSum(Posit32[],Quire).0.num\ := \Posit32::FusedSum(Posit32[],Quire).0.binaryOperationResult.1\;
                            
                            if (\Posit32::FusedSum(Posit32[],Quire).0._State\ = \Posit32::FusedSum(Posit32[],Quire).0._State_14\) then 
                                \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_8\;
                            end if;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Quire Posit32::op_Explicit(Posit32).0._StateMachine\: process (\Clock\) 
        Variable \Quire Posit32::op_Explicit(Posit32).0._State\: \Quire Posit32::op_Explicit(Posit32).0._States\ := \Quire Posit32::op_Explicit(Posit32).0._State_0\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.x\: \Lombiq.Arithmetics.Posit32\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.array\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
        Variable \Quire Posit32::op_Explicit(Posit32).0.return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.quire\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.return.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.0\: signed(63 downto 0) := to_signed(0, 64);
        Variable \Quire Posit32::op_Explicit(Posit32).0.return.2\: signed(15 downto 0) := to_signed(0, 16);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.return.3\: \Lombiq.Arithmetics.Quire\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Quire Posit32::op_Explicit(Posit32).0._Finished\ <= false;
                \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionWithHiddenBit()._Started.0\ <= false;
                \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 64));
                \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= false;
                \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionSize()._Started.0\ <= false;
                \Quire Posit32::op_Explicit(Posit32).0.Posit32::CalculateScaleFactor()._Started.0\ <= false;
                \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\ <= to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ <= false;
                \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_0\;
                \Quire Posit32::op_Explicit(Posit32).0.array\ := (others => to_unsigned(0, 64));
                \Quire Posit32::op_Explicit(Posit32).0.return.0\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.return.1\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.0\ := to_signed(0, 64);
                \Quire Posit32::op_Explicit(Posit32).0.return.2\ := to_signed(0, 16);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.1\ := to_signed(0, 32);
            else 
                case \Quire Posit32::op_Explicit(Posit32).0._State\ is 
                    when \Quire Posit32::op_Explicit(Posit32).0._State_0\ => 
                        
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._Started\ = true) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_2\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_1\ => 
                        
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._Started\ = true) then 
                            \Quire Posit32::op_Explicit(Posit32).0._Finished\ <= true;
                        else 
                            \Quire Posit32::op_Explicit(Posit32).0._Finished\ <= false;
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_0\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_2\ => 
                        \Quire Posit32::op_Explicit(Posit32).0.x\ := \Quire Posit32::op_Explicit(Posit32).0.x.parameter.In\;
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.array\ := (others => to_unsigned(0, 64));
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionWithHiddenBit().this.parameter.Out.0\ <= \Quire Posit32::op_Explicit(Posit32).0.x\;
                        \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionWithHiddenBit()._Started.0\ <= true;
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_3\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_3\ => 
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionWithHiddenBit()._Started.0\ = \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionWithHiddenBit()._Finished.0\) then 
                            \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionWithHiddenBit()._Started.0\ <= false;
                            \Quire Posit32::op_Explicit(Posit32).0.return.0\ := \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionWithHiddenBit().return.0\;
                            \Quire Posit32::op_Explicit(Posit32).0.array\(to_integer(to_signed(0, 32))) := SmartResize(\Quire Posit32::op_Explicit(Posit32).0.return.0\, 64);
                            
                            
                            
                            
                            
                            
                            
                            \Quire Posit32::op_Explicit(Posit32).0.quire\.\IsNull\ := false;
                            \Quire Posit32::op_Explicit(Posit32).0.quire\.\Size\ := to_unsigned(0, 16);
                            \Quire Posit32::op_Explicit(Posit32).0.quire\.\SegmentCount\ := to_unsigned(0, 16);
                            \Quire Posit32::op_Explicit(Posit32).0.quire\.\Segments\ := (others => to_unsigned(0, 64));
                            
                            
                            \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\ <= \Quire Posit32::op_Explicit(Posit32).0.quire\;
                            \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\ <= \Quire Posit32::op_Explicit(Posit32).0.array\;
                            \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\ <= SmartResize(unsigned(to_signed(0, 32)), 16);
                            \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= true;
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_4\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_4\ => 
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ = \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\) then 
                            \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= false;
                            \Quire Posit32::op_Explicit(Posit32).0.quire\ := \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\;
                            \Quire Posit32::op_Explicit(Posit32).0.array\ := \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\;
                            
                            
                            
                            
                            \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionSize().this.parameter.Out.0\ <= \Quire Posit32::op_Explicit(Posit32).0.x\;
                            \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionSize()._Started.0\ <= true;
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_5\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_5\ => 
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionSize()._Started.0\ = \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionSize()._Finished.0\) then 
                            \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionSize()._Started.0\ <= false;
                            \Quire Posit32::op_Explicit(Posit32).0.return.1\ := \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionSize().return.0\;
                            \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.0\ := to_signed(240, 64) - signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.return.1\), 64));
                            
                            \Quire Posit32::op_Explicit(Posit32).0.Posit32::CalculateScaleFactor().this.parameter.Out.0\ <= \Quire Posit32::op_Explicit(Posit32).0.x\;
                            \Quire Posit32::op_Explicit(Posit32).0.Posit32::CalculateScaleFactor()._Started.0\ <= true;
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_6\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_6\ => 
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0.Posit32::CalculateScaleFactor()._Started.0\ = \Quire Posit32::op_Explicit(Posit32).0.Posit32::CalculateScaleFactor()._Finished.0\) then 
                            \Quire Posit32::op_Explicit(Posit32).0.Posit32::CalculateScaleFactor()._Started.0\ <= false;
                            \Quire Posit32::op_Explicit(Posit32).0.return.2\ := \Quire Posit32::op_Explicit(Posit32).0.Posit32::CalculateScaleFactor().return.0\;
                            \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.1\ := SmartResize(\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.0\ + SmartResize((\Quire Posit32::op_Explicit(Posit32).0.return.2\), 64), 32);
                            
                            \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.Out.0\ <= \Quire Posit32::op_Explicit(Posit32).0.quire\;
                            \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\ <= (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.1\);
                            \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ <= true;
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_7\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_7\ => 
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ = \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\) then 
                            \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ <= false;
                            \Quire Posit32::op_Explicit(Posit32).0.return.3\ := \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).return.0\;
                            \Quire Posit32::op_Explicit(Posit32).0.quire\ := \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.In.0\;
                            \Quire Posit32::op_Explicit(Posit32).0.quire\ := \Quire Posit32::op_Explicit(Posit32).0.return.3\;
                            
                            
                            
                            \Quire Posit32::op_Explicit(Posit32).0.return\ <= \Quire Posit32::op_Explicit(Posit32).0.quire\;
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_1\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Quire::.ctor(UInt64[],UInt16).0._StateMachine\: process (\Clock\) 
        Variable \Quire::.ctor(UInt64[],UInt16).0._State\: \Quire::.ctor(UInt64[],UInt16).0._States\ := \Quire::.ctor(UInt64[],UInt16).0._State_0\;
        Variable \Quire::.ctor(UInt64[],UInt16).0.this\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire::.ctor(UInt64[],UInt16).0.segments\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
        Variable \Quire::.ctor(UInt64[],UInt16).0.size\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire::.ctor(UInt64[],UInt16).0.num\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire::.ctor(UInt64[],UInt16).0.binaryOperationResult.0\: boolean := false;
        Variable \Quire::.ctor(UInt64[],UInt16).0.binaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Quire::.ctor(UInt64[],UInt16).0._Finished\ <= false;
                \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.Out\ <= (others => to_unsigned(0, 64));
                \Quire::.ctor(UInt64[],UInt16).0._State\ := \Quire::.ctor(UInt64[],UInt16).0._State_0\;
                \Quire::.ctor(UInt64[],UInt16).0.segments\ := (others => to_unsigned(0, 64));
                \Quire::.ctor(UInt64[],UInt16).0.size\ := to_unsigned(0, 16);
                \Quire::.ctor(UInt64[],UInt16).0.num\ := to_signed(0, 32);
                \Quire::.ctor(UInt64[],UInt16).0.binaryOperationResult.0\ := false;
                \Quire::.ctor(UInt64[],UInt16).0.binaryOperationResult.1\ := to_signed(0, 32);
            else 
                case \Quire::.ctor(UInt64[],UInt16).0._State\ is 
                    when \Quire::.ctor(UInt64[],UInt16).0._State_0\ => 
                        
                        
                        if (\Quire::.ctor(UInt64[],UInt16).0._Started\ = true) then 
                            \Quire::.ctor(UInt64[],UInt16).0._State\ := \Quire::.ctor(UInt64[],UInt16).0._State_2\;
                        end if;
                        
                    when \Quire::.ctor(UInt64[],UInt16).0._State_1\ => 
                        
                        
                        if (\Quire::.ctor(UInt64[],UInt16).0._Started\ = true) then 
                            \Quire::.ctor(UInt64[],UInt16).0._Finished\ <= true;
                        else 
                            \Quire::.ctor(UInt64[],UInt16).0._Finished\ <= false;
                            \Quire::.ctor(UInt64[],UInt16).0._State\ := \Quire::.ctor(UInt64[],UInt16).0._State_0\;
                        end if;
                        
                        \Quire::.ctor(UInt64[],UInt16).0.this.parameter.Out\ <= \Quire::.ctor(UInt64[],UInt16).0.this\;
                        \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.Out\ <= \Quire::.ctor(UInt64[],UInt16).0.segments\;
                        
                    when \Quire::.ctor(UInt64[],UInt16).0._State_2\ => 
                        \Quire::.ctor(UInt64[],UInt16).0.this\ := \Quire::.ctor(UInt64[],UInt16).0.this.parameter.In\;
                        \Quire::.ctor(UInt64[],UInt16).0.segments\ := \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.In\;
                        \Quire::.ctor(UInt64[],UInt16).0.size\ := \Quire::.ctor(UInt64[],UInt16).0.size.parameter.In\;
                        
                        
                        
                        \Quire::.ctor(UInt64[],UInt16).0.this\.\SegmentCount\ := to_unsigned(8, 16);
                        
                        
                        
                        \Quire::.ctor(UInt64[],UInt16).0.this\.\Size\ := SmartResize(unsigned(to_signed(0, 32)), 16);
                        
                        
                        
                        \Quire::.ctor(UInt64[],UInt16).0.this\.\Segments\ := (others => to_unsigned(0, 64));
                        
                        
                        
                        \Quire::.ctor(UInt64[],UInt16).0.this\.\Segments\ := \Quire::.ctor(UInt64[],UInt16).0.segments\(0 to 7);
                        
                        
                        
                        
                        
                        
                        \Quire::.ctor(UInt64[],UInt16).0.num\ := to_signed(8, 32);
                        
                        
                        
                        
                        
                        
                        
                        \Quire::.ctor(UInt64[],UInt16).0._State\ := \Quire::.ctor(UInt64[],UInt16).0._State_3\;
                        
                    when \Quire::.ctor(UInt64[],UInt16).0._State_3\ => 
                        
                        
                        \Quire::.ctor(UInt64[],UInt16).0.binaryOperationResult.0\ := (\Quire::.ctor(UInt64[],UInt16).0.num\) < to_signed(8, 32);
                        if (\Quire::.ctor(UInt64[],UInt16).0.binaryOperationResult.0\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire::.ctor(UInt64[],UInt16).0.this\.\Segments\(to_integer(\Quire::.ctor(UInt64[],UInt16).0.num\)) := to_unsigned(0, 64);
                            
                            
                            
                            \Quire::.ctor(UInt64[],UInt16).0.binaryOperationResult.1\ := \Quire::.ctor(UInt64[],UInt16).0.num\ + to_signed(1, 32);
                            \Quire::.ctor(UInt64[],UInt16).0.num\ := \Quire::.ctor(UInt64[],UInt16).0.binaryOperationResult.1\;
                        else 
                            \Quire::.ctor(UInt64[],UInt16).0._State\ := \Quire::.ctor(UInt64[],UInt16).0._State_4\;
                        end if;
                        
                    when \Quire::.ctor(UInt64[],UInt16).0._State_4\ => 
                        
                        \Quire::.ctor(UInt64[],UInt16).0._State\ := \Quire::.ctor(UInt64[],UInt16).0._State_1\;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Quire::.ctor(UInt32,UInt16).0._StateMachine\: process (\Clock\) 
        Variable \Quire::.ctor(UInt32,UInt16).0._State\: \Quire::.ctor(UInt32,UInt16).0._States\ := \Quire::.ctor(UInt32,UInt16).0._State_0\;
        Variable \Quire::.ctor(UInt32,UInt16).0.this\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire::.ctor(UInt32,UInt16).0.firstSegment\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire::.ctor(UInt32,UInt16).0.size\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire::.ctor(UInt32,UInt16).0.conditional508ca86de85a5da84bb49b246fc4b145e1352a0547a47e41f17ab54c68695517\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire::.ctor(UInt32,UInt16).0.remainderOperand0c439d9dfdc1e321f9179f8d0530a346aae5aa4d433af564a6e961f787b90b5b\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.3\: boolean := false;
        Variable \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.4\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.5\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire::.ctor(UInt32,UInt16).0.num\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.6\: boolean := false;
        Variable \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.7\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Quire::.ctor(UInt32,UInt16).0._Finished\ <= false;
                \Quire::.ctor(UInt32,UInt16).0._State\ := \Quire::.ctor(UInt32,UInt16).0._State_0\;
                \Quire::.ctor(UInt32,UInt16).0.firstSegment\ := to_unsigned(0, 32);
                \Quire::.ctor(UInt32,UInt16).0.size\ := to_unsigned(0, 16);
                \Quire::.ctor(UInt32,UInt16).0.conditional508ca86de85a5da84bb49b246fc4b145e1352a0547a47e41f17ab54c68695517\ := to_signed(0, 32);
                \Quire::.ctor(UInt32,UInt16).0.remainderOperand0c439d9dfdc1e321f9179f8d0530a346aae5aa4d433af564a6e961f787b90b5b\ := to_signed(0, 32);
                \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.0\ := to_signed(0, 32);
                \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.1\ := to_signed(0, 32);
                \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.2\ := to_signed(0, 32);
                \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.3\ := false;
                \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.4\ := to_signed(0, 32);
                \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.5\ := to_unsigned(0, 16);
                \Quire::.ctor(UInt32,UInt16).0.num\ := to_signed(0, 32);
                \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.6\ := false;
                \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.7\ := to_signed(0, 32);
            else 
                case \Quire::.ctor(UInt32,UInt16).0._State\ is 
                    when \Quire::.ctor(UInt32,UInt16).0._State_0\ => 
                        
                        
                        if (\Quire::.ctor(UInt32,UInt16).0._Started\ = true) then 
                            \Quire::.ctor(UInt32,UInt16).0._State\ := \Quire::.ctor(UInt32,UInt16).0._State_2\;
                        end if;
                        
                    when \Quire::.ctor(UInt32,UInt16).0._State_1\ => 
                        
                        
                        if (\Quire::.ctor(UInt32,UInt16).0._Started\ = true) then 
                            \Quire::.ctor(UInt32,UInt16).0._Finished\ <= true;
                        else 
                            \Quire::.ctor(UInt32,UInt16).0._Finished\ <= false;
                            \Quire::.ctor(UInt32,UInt16).0._State\ := \Quire::.ctor(UInt32,UInt16).0._State_0\;
                        end if;
                        
                        \Quire::.ctor(UInt32,UInt16).0.this.parameter.Out\ <= \Quire::.ctor(UInt32,UInt16).0.this\;
                        
                    when \Quire::.ctor(UInt32,UInt16).0._State_2\ => 
                        \Quire::.ctor(UInt32,UInt16).0.this\ := \Quire::.ctor(UInt32,UInt16).0.this.parameter.In\;
                        \Quire::.ctor(UInt32,UInt16).0.firstSegment\ := \Quire::.ctor(UInt32,UInt16).0.firstSegment.parameter.In\;
                        \Quire::.ctor(UInt32,UInt16).0.size\ := \Quire::.ctor(UInt32,UInt16).0.size.parameter.In\;
                        
                        
                        
                        \Quire::.ctor(UInt32,UInt16).0.this\.\Size\ := \Quire::.ctor(UInt32,UInt16).0.size\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire::.ctor(UInt32,UInt16).0.remainderOperand0c439d9dfdc1e321f9179f8d0530a346aae5aa4d433af564a6e961f787b90b5b\ := signed(SmartResize(\Quire::.ctor(UInt32,UInt16).0.size\, 32));
                        
                        
                        
                        
                        
                        
                        
                        \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.0\ := \Quire::.ctor(UInt32,UInt16).0.remainderOperand0c439d9dfdc1e321f9179f8d0530a346aae5aa4d433af564a6e961f787b90b5b\ / to_signed(32, 32);
                        \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.1\ := SmartResize(\Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.0\ * to_signed(32, 32), 32);
                        \Quire::.ctor(UInt32,UInt16).0._State\ := \Quire::.ctor(UInt32,UInt16).0._State_3\;
                        
                    when \Quire::.ctor(UInt32,UInt16).0._State_3\ => 
                        
                        \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.2\ := \Quire::.ctor(UInt32,UInt16).0.remainderOperand0c439d9dfdc1e321f9179f8d0530a346aae5aa4d433af564a6e961f787b90b5b\ - \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.1\;
                        \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.3\ := \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.2\ /= to_signed(0, 32);

                        
                        
                        
                        

                        if ((\Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.3\)) then 
                            \Quire::.ctor(UInt32,UInt16).0._State\ := \Quire::.ctor(UInt32,UInt16).0._State_5\;
                        else 
                            \Quire::.ctor(UInt32,UInt16).0._State\ := \Quire::.ctor(UInt32,UInt16).0._State_6\;
                        end if;
                        
                    when \Quire::.ctor(UInt32,UInt16).0._State_4\ => 
                        
                        
                        
                        
                        \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.4\ := shift_right(signed(SmartResize((\Quire::.ctor(UInt32,UInt16).0.size\), 32)), to_integer(unsigned(SmartResize(to_signed(6, 32), 5) and "11111")));
                        \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.5\ := SmartResize(unsigned((\Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.4\) + (\Quire::.ctor(UInt32,UInt16).0.conditional508ca86de85a5da84bb49b246fc4b145e1352a0547a47e41f17ab54c68695517\)), 16);
                        \Quire::.ctor(UInt32,UInt16).0.this\.\SegmentCount\ := (\Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.5\);
                        
                        
                        
                        \Quire::.ctor(UInt32,UInt16).0.this\.\Segments\ := (others => to_unsigned(0, 64));
                        
                        
                        
                        \Quire::.ctor(UInt32,UInt16).0.this\.\Segments\(to_integer(to_signed(0, 32))) := SmartResize(to_unsigned(1, 32), 64);
                        
                        
                        
                        
                        
                        
                        \Quire::.ctor(UInt32,UInt16).0.num\ := to_signed(1, 32);
                        
                        
                        
                        
                        
                        
                        
                        \Quire::.ctor(UInt32,UInt16).0._State\ := \Quire::.ctor(UInt32,UInt16).0._State_7\;
                        
                    when \Quire::.ctor(UInt32,UInt16).0._State_5\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire::.ctor(UInt32,UInt16).0.conditional508ca86de85a5da84bb49b246fc4b145e1352a0547a47e41f17ab54c68695517\ := to_signed(1, 32);
                        
                        if (\Quire::.ctor(UInt32,UInt16).0._State\ = \Quire::.ctor(UInt32,UInt16).0._State_5\) then 
                            \Quire::.ctor(UInt32,UInt16).0._State\ := \Quire::.ctor(UInt32,UInt16).0._State_4\;
                        end if;
                        
                    when \Quire::.ctor(UInt32,UInt16).0._State_6\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire::.ctor(UInt32,UInt16).0.conditional508ca86de85a5da84bb49b246fc4b145e1352a0547a47e41f17ab54c68695517\ := to_signed(0, 32);
                        
                        if (\Quire::.ctor(UInt32,UInt16).0._State\ = \Quire::.ctor(UInt32,UInt16).0._State_6\) then 
                            \Quire::.ctor(UInt32,UInt16).0._State\ := \Quire::.ctor(UInt32,UInt16).0._State_4\;
                        end if;
                        
                    when \Quire::.ctor(UInt32,UInt16).0._State_7\ => 
                        
                        
                        \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.6\ := (\Quire::.ctor(UInt32,UInt16).0.num\) < signed(SmartResize((\Quire::.ctor(UInt32,UInt16).0.this\.\SegmentCount\), 32));
                        if (\Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.6\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire::.ctor(UInt32,UInt16).0.this\.\Segments\(to_integer(\Quire::.ctor(UInt32,UInt16).0.num\)) := to_unsigned(0, 64);
                            
                            
                            
                            \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.7\ := \Quire::.ctor(UInt32,UInt16).0.num\ + to_signed(1, 32);
                            \Quire::.ctor(UInt32,UInt16).0.num\ := \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.7\;
                        else 
                            \Quire::.ctor(UInt32,UInt16).0._State\ := \Quire::.ctor(UInt32,UInt16).0._State_8\;
                        end if;
                        
                    when \Quire::.ctor(UInt32,UInt16).0._State_8\ => 
                        
                        \Quire::.ctor(UInt32,UInt16).0._State\ := \Quire::.ctor(UInt32,UInt16).0._State_1\;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Quire Quire::op_Addition(Quire,Quire).0._StateMachine\: process (\Clock\) 
        Variable \Quire Quire::op_Addition(Quire,Quire).0._State\: \Quire Quire::op_Addition(Quire,Quire).0._States\ := \Quire Quire::op_Addition(Quire,Quire).0._State_0\;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.left\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.right\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.0\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.1\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.2\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.array\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
        Variable \Quire Quire::op_Addition(Quire,Quire).0.flag\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.num\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.num2\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.num3\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.3\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.4\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.flag2\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.5\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.6\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.7\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.flag3\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.8\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.9\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.10\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.b\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.conditional746a1c636f616ff3623be4e48942688719382078a087cbdab0e2c998303da9ba\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.conditionalc042a0f1121d35344a49419953dc5f52591ee75c13d7b4714794eeff7d14bf49\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.conditionalae2b32de30beca2038d02dc985eb3cd14f87df2ffaa1520711b83d6b5e0acd70\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.11\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.12\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.13\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.14\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.15\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.16\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.17\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.18\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.19\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.20\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.21\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.22\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.23\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.objectd7f66d6090a3f51dbf9c6b85d3744cbaf909687ec9d3f52027672e9a5e2ece9d\: \Lombiq.Arithmetics.Quire\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Quire Quire::op_Addition(Quire,Quire).0._Finished\ <= false;
                \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 64));
                \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= false;
                \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_0\;
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.0\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.1\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.2\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.array\ := (others => to_unsigned(0, 64));
                \Quire Quire::op_Addition(Quire,Quire).0.flag\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.num\ := to_unsigned(0, 16);
                \Quire Quire::op_Addition(Quire,Quire).0.num2\ := to_unsigned(0, 16);
                \Quire Quire::op_Addition(Quire,Quire).0.num3\ := to_unsigned(0, 16);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.3\ := to_signed(0, 32);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.4\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.flag2\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.5\ := to_unsigned(0, 64);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.6\ := to_unsigned(0, 64);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.7\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.flag3\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.8\ := to_unsigned(0, 64);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.9\ := to_unsigned(0, 64);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.10\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.b\ := to_unsigned(0, 8);
                \Quire Quire::op_Addition(Quire,Quire).0.conditional746a1c636f616ff3623be4e48942688719382078a087cbdab0e2c998303da9ba\ := to_signed(0, 32);
                \Quire Quire::op_Addition(Quire,Quire).0.conditionalc042a0f1121d35344a49419953dc5f52591ee75c13d7b4714794eeff7d14bf49\ := to_signed(0, 32);
                \Quire Quire::op_Addition(Quire,Quire).0.conditionalae2b32de30beca2038d02dc985eb3cd14f87df2ffaa1520711b83d6b5e0acd70\ := to_signed(0, 32);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.11\ := to_signed(0, 32);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.12\ := to_unsigned(0, 8);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.13\ := to_signed(0, 32);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.14\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.15\ := to_unsigned(0, 64);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.16\ := to_unsigned(0, 64);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.17\ := to_signed(0, 32);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.18\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.19\ := to_unsigned(0, 16);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.20\ := to_signed(0, 32);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.21\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.22\ := to_unsigned(0, 16);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.23\ := to_unsigned(0, 16);
            else 
                case \Quire Quire::op_Addition(Quire,Quire).0._State\ is 
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_0\ => 
                        
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._Started\ = true) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_2\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_1\ => 
                        
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._Started\ = true) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._Finished\ <= true;
                        else 
                            \Quire Quire::op_Addition(Quire,Quire).0._Finished\ <= false;
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_0\;
                        end if;
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.left.parameter.Out\ <= \Quire Quire::op_Addition(Quire,Quire).0.left\;
                        \Quire Quire::op_Addition(Quire,Quire).0.right.parameter.Out\ <= \Quire Quire::op_Addition(Quire,Quire).0.right\;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_2\ => 
                        \Quire Quire::op_Addition(Quire,Quire).0.left\ := \Quire Quire::op_Addition(Quire,Quire).0.left.parameter.In\;
                        \Quire Quire::op_Addition(Quire,Quire).0.right\ := \Quire Quire::op_Addition(Quire,Quire).0.right.parameter.In\;
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.0\ := signed(SmartResize((\Quire Quire::op_Addition(Quire,Quire).0.left\.\SegmentCount\), 32)) = to_signed(0, 32);
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.1\ := signed(SmartResize((\Quire Quire::op_Addition(Quire,Quire).0.right\.\SegmentCount\), 32)) = to_signed(0, 32);
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.2\ := \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.0\ or \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.1\;

                        
                        
                        

                        if (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.2\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_4\;
                        else 
                            
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_3\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_3\ => 
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.array\ := (others => to_unsigned(0, 64));
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.flag\ := false;
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.num\ := SmartResize(unsigned(to_signed(0, 32)), 16);
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.num2\ := SmartResize(unsigned(to_signed(0, 32)), 16);
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.num3\ := SmartResize(unsigned(to_signed(0, 32)), 16);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_5\;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_4\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.return\ <= \Quire Quire::op_Addition(Quire,Quire).0.left\;
                        \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_1\;
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._State\ = \Quire Quire::op_Addition(Quire,Quire).0._State_4\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_3\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_5\ => 
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.3\ := shift_left(signed(SmartResize((\Quire Quire::op_Addition(Quire,Quire).0.left\.\SegmentCount\), 32)), to_integer(unsigned(SmartResize(to_signed(6, 32), 5))));
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.4\ := signed(SmartResize((\Quire Quire::op_Addition(Quire,Quire).0.num3\), 32)) < (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.3\);
                        if (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.4\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_7\;
                        else 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_6\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_6\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.objectd7f66d6090a3f51dbf9c6b85d3744cbaf909687ec9d3f52027672e9a5e2ece9d\.\IsNull\ := false;
                        \Quire Quire::op_Addition(Quire,Quire).0.objectd7f66d6090a3f51dbf9c6b85d3744cbaf909687ec9d3f52027672e9a5e2ece9d\.\Size\ := to_unsigned(0, 16);
                        \Quire Quire::op_Addition(Quire,Quire).0.objectd7f66d6090a3f51dbf9c6b85d3744cbaf909687ec9d3f52027672e9a5e2ece9d\.\SegmentCount\ := to_unsigned(0, 16);
                        \Quire Quire::op_Addition(Quire,Quire).0.objectd7f66d6090a3f51dbf9c6b85d3744cbaf909687ec9d3f52027672e9a5e2ece9d\.\Segments\ := (others => to_unsigned(0, 64));
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\ <= \Quire Quire::op_Addition(Quire,Quire).0.objectd7f66d6090a3f51dbf9c6b85d3744cbaf909687ec9d3f52027672e9a5e2ece9d\;
                        \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\ <= \Quire Quire::op_Addition(Quire,Quire).0.array\;
                        \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\ <= SmartResize(unsigned(to_signed(0, 32)), 16);
                        \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= true;
                        \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_28\;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_7\ => 
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.5\ := SmartResize(shift_right(\Quire Quire::op_Addition(Quire,Quire).0.left\.\Segments\(to_integer(\Quire Quire::op_Addition(Quire,Quire).0.num\)), to_integer(unsigned(SmartResize(signed(SmartResize(\Quire Quire::op_Addition(Quire,Quire).0.num2\, 32)), 6) and "111111"))), 64);
                        \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_8\;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_8\ => 
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.6\ := (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.5\) and to_unsigned(1, 64);
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.7\ := (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.6\) = to_unsigned(1, 64);
                        \Quire Quire::op_Addition(Quire,Quire).0.flag2\ := \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.7\;
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_9\;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_9\ => 
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.8\ := SmartResize(shift_right(\Quire Quire::op_Addition(Quire,Quire).0.right\.\Segments\(to_integer(\Quire Quire::op_Addition(Quire,Quire).0.num\)), to_integer(unsigned(SmartResize(signed(SmartResize(\Quire Quire::op_Addition(Quire,Quire).0.num2\, 32)), 6) and "111111"))), 64);
                        \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_10\;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_10\ => 
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.9\ := (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.8\) and to_unsigned(1, 64);
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.10\ := (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.9\) = to_unsigned(1, 64);
                        \Quire Quire::op_Addition(Quire,Quire).0.flag3\ := \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.10\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        

                        
                        
                        
                        

                        if (\Quire Quire::op_Addition(Quire,Quire).0.flag2\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_12\;
                        else 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_13\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_11\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        

                        
                        
                        
                        

                        if (\Quire Quire::op_Addition(Quire,Quire).0.flag3\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_15\;
                        else 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_16\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_12\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.conditional746a1c636f616ff3623be4e48942688719382078a087cbdab0e2c998303da9ba\ := to_signed(1, 32);
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._State\ = \Quire Quire::op_Addition(Quire,Quire).0._State_12\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_11\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_13\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.conditional746a1c636f616ff3623be4e48942688719382078a087cbdab0e2c998303da9ba\ := to_signed(0, 32);
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._State\ = \Quire Quire::op_Addition(Quire,Quire).0._State_13\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_11\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_14\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        

                        
                        
                        
                        

                        if (\Quire Quire::op_Addition(Quire,Quire).0.flag\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_18\;
                        else 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_19\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_15\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.conditionalc042a0f1121d35344a49419953dc5f52591ee75c13d7b4714794eeff7d14bf49\ := to_signed(1, 32);
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._State\ = \Quire Quire::op_Addition(Quire,Quire).0._State_15\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_14\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_16\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.conditionalc042a0f1121d35344a49419953dc5f52591ee75c13d7b4714794eeff7d14bf49\ := to_signed(0, 32);
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._State\ = \Quire Quire::op_Addition(Quire,Quire).0._State_16\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_14\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_17\ => 
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.11\ := (\Quire Quire::op_Addition(Quire,Quire).0.conditional746a1c636f616ff3623be4e48942688719382078a087cbdab0e2c998303da9ba\) + (\Quire Quire::op_Addition(Quire,Quire).0.conditionalc042a0f1121d35344a49419953dc5f52591ee75c13d7b4714794eeff7d14bf49\);
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.12\ := SmartResize(unsigned(\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.11\ + (\Quire Quire::op_Addition(Quire,Quire).0.conditionalae2b32de30beca2038d02dc985eb3cd14f87df2ffaa1520711b83d6b5e0acd70\)), 8);
                        \Quire Quire::op_Addition(Quire,Quire).0.b\ := (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.12\);
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.13\ := signed(SmartResize((\Quire Quire::op_Addition(Quire,Quire).0.b\), 32)) and to_signed(1, 32);
                        \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_20\;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_18\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.conditionalae2b32de30beca2038d02dc985eb3cd14f87df2ffaa1520711b83d6b5e0acd70\ := to_signed(1, 32);
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._State\ = \Quire Quire::op_Addition(Quire,Quire).0._State_18\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_17\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_19\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.conditionalae2b32de30beca2038d02dc985eb3cd14f87df2ffaa1520711b83d6b5e0acd70\ := to_signed(0, 32);
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._State\ = \Quire Quire::op_Addition(Quire,Quire).0._State_19\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_17\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_20\ => 
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.14\ := (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.13\) = to_signed(1, 32);

                        
                        
                        

                        if (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.14\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_22\;
                        else 
                            
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_21\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_21\ => 
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.17\ := shift_right(signed(SmartResize((\Quire Quire::op_Addition(Quire,Quire).0.b\), 32)), to_integer(unsigned(SmartResize(to_signed(1, 32), 5) and "11111")));
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.18\ := \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.17\ = to_signed(1, 32);
                        \Quire Quire::op_Addition(Quire,Quire).0.flag\ := \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.18\;
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_24\;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_22\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.15\ := SmartResize(unsigned(shift_left(to_signed(1, 64), to_integer(unsigned(SmartResize(signed(SmartResize(\Quire Quire::op_Addition(Quire,Quire).0.num2\, 32)), 6))))), 64);
                        \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_23\;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_23\ => 
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.16\ := \Quire Quire::op_Addition(Quire,Quire).0.array\(to_integer(\Quire Quire::op_Addition(Quire,Quire).0.num\)) + (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.15\);
                        \Quire Quire::op_Addition(Quire,Quire).0.array\(to_integer(\Quire Quire::op_Addition(Quire,Quire).0.num\)) := \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.16\;
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._State\ = \Quire Quire::op_Addition(Quire,Quire).0._State_23\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_21\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_24\ => 
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.19\ := SmartResize(unsigned(signed(SmartResize((\Quire Quire::op_Addition(Quire,Quire).0.num2\), 32)) + to_signed(1, 32)), 16);
                        \Quire Quire::op_Addition(Quire,Quire).0.num2\ := (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.19\);
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.20\ := shift_right(signed(SmartResize((\Quire Quire::op_Addition(Quire,Quire).0.num2\), 32)), to_integer(unsigned(SmartResize(to_signed(6, 32), 5) and "11111")));
                        \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_25\;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_25\ => 
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.21\ := \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.20\ = to_signed(1, 32);

                        
                        
                        

                        if (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.21\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_27\;
                        else 
                            
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_26\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_26\ => 
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.23\ := SmartResize(unsigned(signed(SmartResize((\Quire Quire::op_Addition(Quire,Quire).0.num3\), 32)) + to_signed(1, 32)), 16);
                        \Quire Quire::op_Addition(Quire,Quire).0.num3\ := (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.23\);
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._State\ = \Quire Quire::op_Addition(Quire,Quire).0._State_26\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_5\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_27\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.num2\ := SmartResize(unsigned(to_signed(0, 32)), 16);
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.22\ := SmartResize(unsigned(signed(SmartResize((\Quire Quire::op_Addition(Quire,Quire).0.num\), 32)) + to_signed(1, 32)), 16);
                        \Quire Quire::op_Addition(Quire,Quire).0.num\ := (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.22\);
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._State\ = \Quire Quire::op_Addition(Quire,Quire).0._State_27\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_26\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_28\ => 
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ = \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= false;
                            \Quire Quire::op_Addition(Quire,Quire).0.objectd7f66d6090a3f51dbf9c6b85d3744cbaf909687ec9d3f52027672e9a5e2ece9d\ := \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\;
                            \Quire Quire::op_Addition(Quire,Quire).0.array\ := \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\;
                            
                            
                            
                            \Quire Quire::op_Addition(Quire,Quire).0.return\ <= \Quire Quire::op_Addition(Quire,Quire).0.objectd7f66d6090a3f51dbf9c6b85d3744cbaf909687ec9d3f52027672e9a5e2ece9d\;
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_1\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Quire Quire::op_Addition(Quire,UInt32).0._StateMachine\: process (\Clock\) 
        Variable \Quire Quire::op_Addition(Quire,UInt32).0._State\: \Quire Quire::op_Addition(Quire,UInt32).0._States\ := \Quire Quire::op_Addition(Quire,UInt32).0._State_0\;
        Variable \Quire Quire::op_Addition(Quire,UInt32).0.left\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire Quire::op_Addition(Quire,UInt32).0.right\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Quire::op_Addition(Quire,UInt32).0.object2b25f3fa9b50e7492d78b34e15a583b8300db89f75b5c7cb2910bbab85a19ff0\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire Quire::op_Addition(Quire,UInt32).0.binaryOperationResult.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_Addition(Quire,UInt32).0.return.0\: \Lombiq.Arithmetics.Quire\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Quire Quire::op_Addition(Quire,UInt32).0._Finished\ <= false;
                \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).firstSegment.parameter.Out.0\ <= to_unsigned(0, 32);
                \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Started.0\ <= false;
                \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\ <= false;
                \Quire Quire::op_Addition(Quire,UInt32).0._State\ := \Quire Quire::op_Addition(Quire,UInt32).0._State_0\;
                \Quire Quire::op_Addition(Quire,UInt32).0.right\ := to_unsigned(0, 32);
                \Quire Quire::op_Addition(Quire,UInt32).0.binaryOperationResult.0\ := to_unsigned(0, 16);
            else 
                case \Quire Quire::op_Addition(Quire,UInt32).0._State\ is 
                    when \Quire Quire::op_Addition(Quire,UInt32).0._State_0\ => 
                        
                        
                        if (\Quire Quire::op_Addition(Quire,UInt32).0._Started\ = true) then 
                            \Quire Quire::op_Addition(Quire,UInt32).0._State\ := \Quire Quire::op_Addition(Quire,UInt32).0._State_2\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,UInt32).0._State_1\ => 
                        
                        
                        if (\Quire Quire::op_Addition(Quire,UInt32).0._Started\ = true) then 
                            \Quire Quire::op_Addition(Quire,UInt32).0._Finished\ <= true;
                        else 
                            \Quire Quire::op_Addition(Quire,UInt32).0._Finished\ <= false;
                            \Quire Quire::op_Addition(Quire,UInt32).0._State\ := \Quire Quire::op_Addition(Quire,UInt32).0._State_0\;
                        end if;
                        
                        \Quire Quire::op_Addition(Quire,UInt32).0.left.parameter.Out\ <= \Quire Quire::op_Addition(Quire,UInt32).0.left\;
                        
                    when \Quire Quire::op_Addition(Quire,UInt32).0._State_2\ => 
                        \Quire Quire::op_Addition(Quire,UInt32).0.left\ := \Quire Quire::op_Addition(Quire,UInt32).0.left.parameter.In\;
                        \Quire Quire::op_Addition(Quire,UInt32).0.right\ := \Quire Quire::op_Addition(Quire,UInt32).0.right.parameter.In\;
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,UInt32).0.object2b25f3fa9b50e7492d78b34e15a583b8300db89f75b5c7cb2910bbab85a19ff0\.\IsNull\ := false;
                        \Quire Quire::op_Addition(Quire,UInt32).0.object2b25f3fa9b50e7492d78b34e15a583b8300db89f75b5c7cb2910bbab85a19ff0\.\Size\ := to_unsigned(0, 16);
                        \Quire Quire::op_Addition(Quire,UInt32).0.object2b25f3fa9b50e7492d78b34e15a583b8300db89f75b5c7cb2910bbab85a19ff0\.\SegmentCount\ := to_unsigned(0, 16);
                        \Quire Quire::op_Addition(Quire,UInt32).0.object2b25f3fa9b50e7492d78b34e15a583b8300db89f75b5c7cb2910bbab85a19ff0\.\Segments\ := (others => to_unsigned(0, 64));
                        
                        \Quire Quire::op_Addition(Quire,UInt32).0.binaryOperationResult.0\ := SmartResize(unsigned(shift_left(signed(SmartResize((\Quire Quire::op_Addition(Quire,UInt32).0.left\.\SegmentCount\), 32)), to_integer(unsigned(SmartResize(to_signed(6, 32), 5))))), 16);
                        
                        \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).this.parameter.Out.0\ <= \Quire Quire::op_Addition(Quire,UInt32).0.object2b25f3fa9b50e7492d78b34e15a583b8300db89f75b5c7cb2910bbab85a19ff0\;
                        \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).firstSegment.parameter.Out.0\ <= to_unsigned(1, 32);
                        \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).size.parameter.Out.0\ <= (\Quire Quire::op_Addition(Quire,UInt32).0.binaryOperationResult.0\);
                        \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Started.0\ <= true;
                        \Quire Quire::op_Addition(Quire,UInt32).0._State\ := \Quire Quire::op_Addition(Quire,UInt32).0._State_3\;
                        
                    when \Quire Quire::op_Addition(Quire,UInt32).0._State_3\ => 
                        
                        if (\Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Started.0\ = \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Finished.0\) then 
                            \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Started.0\ <= false;
                            \Quire Quire::op_Addition(Quire,UInt32).0.object2b25f3fa9b50e7492d78b34e15a583b8300db89f75b5c7cb2910bbab85a19ff0\ := \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).this.parameter.In.0\;
                            
                            
                            
                            
                            \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.Out.0\ <= \Quire Quire::op_Addition(Quire,UInt32).0.left\;
                            \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.Out.0\ <= \Quire Quire::op_Addition(Quire,UInt32).0.object2b25f3fa9b50e7492d78b34e15a583b8300db89f75b5c7cb2910bbab85a19ff0\;
                            \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\ <= true;
                            \Quire Quire::op_Addition(Quire,UInt32).0._State\ := \Quire Quire::op_Addition(Quire,UInt32).0._State_4\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,UInt32).0._State_4\ => 
                        
                        if (\Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\ = \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\) then 
                            \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\ <= false;
                            \Quire Quire::op_Addition(Quire,UInt32).0.return.0\ := \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).return.0\;
                            \Quire Quire::op_Addition(Quire,UInt32).0.left\ := \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.In.0\;
                            \Quire Quire::op_Addition(Quire,UInt32).0.object2b25f3fa9b50e7492d78b34e15a583b8300db89f75b5c7cb2910bbab85a19ff0\ := \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.In.0\;
                            \Quire Quire::op_Addition(Quire,UInt32).0.return\ <= \Quire Quire::op_Addition(Quire,UInt32).0.return.0\;
                            \Quire Quire::op_Addition(Quire,UInt32).0._State\ := \Quire Quire::op_Addition(Quire,UInt32).0._State_1\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Quire Quire::op_OnesComplement(Quire).0._StateMachine\: process (\Clock\) 
        Variable \Quire Quire::op_OnesComplement(Quire).0._State\: \Quire Quire::op_OnesComplement(Quire).0._States\ := \Quire Quire::op_OnesComplement(Quire).0._State_0\;
        Variable \Quire Quire::op_OnesComplement(Quire).0.q\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire Quire::op_OnesComplement(Quire).0.num\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_OnesComplement(Quire).0.binaryOperationResult.0\: boolean := false;
        Variable \Quire Quire::op_OnesComplement(Quire).0.unaryOperationResult.0\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_OnesComplement(Quire).0.binaryOperationResult.1\: unsigned(15 downto 0) := to_unsigned(0, 16);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Quire Quire::op_OnesComplement(Quire).0._Finished\ <= false;
                \Quire Quire::op_OnesComplement(Quire).0._State\ := \Quire Quire::op_OnesComplement(Quire).0._State_0\;
                \Quire Quire::op_OnesComplement(Quire).0.num\ := to_unsigned(0, 16);
                \Quire Quire::op_OnesComplement(Quire).0.binaryOperationResult.0\ := false;
                \Quire Quire::op_OnesComplement(Quire).0.unaryOperationResult.0\ := to_unsigned(0, 64);
                \Quire Quire::op_OnesComplement(Quire).0.binaryOperationResult.1\ := to_unsigned(0, 16);
            else 
                case \Quire Quire::op_OnesComplement(Quire).0._State\ is 
                    when \Quire Quire::op_OnesComplement(Quire).0._State_0\ => 
                        
                        
                        if (\Quire Quire::op_OnesComplement(Quire).0._Started\ = true) then 
                            \Quire Quire::op_OnesComplement(Quire).0._State\ := \Quire Quire::op_OnesComplement(Quire).0._State_2\;
                        end if;
                        
                    when \Quire Quire::op_OnesComplement(Quire).0._State_1\ => 
                        
                        
                        if (\Quire Quire::op_OnesComplement(Quire).0._Started\ = true) then 
                            \Quire Quire::op_OnesComplement(Quire).0._Finished\ <= true;
                        else 
                            \Quire Quire::op_OnesComplement(Quire).0._Finished\ <= false;
                            \Quire Quire::op_OnesComplement(Quire).0._State\ := \Quire Quire::op_OnesComplement(Quire).0._State_0\;
                        end if;
                        
                        \Quire Quire::op_OnesComplement(Quire).0.q.parameter.Out\ <= \Quire Quire::op_OnesComplement(Quire).0.q\;
                        
                    when \Quire Quire::op_OnesComplement(Quire).0._State_2\ => 
                        \Quire Quire::op_OnesComplement(Quire).0.q\ := \Quire Quire::op_OnesComplement(Quire).0.q.parameter.In\;
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_OnesComplement(Quire).0.num\ := SmartResize(unsigned(to_signed(0, 32)), 16);
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_OnesComplement(Quire).0._State\ := \Quire Quire::op_OnesComplement(Quire).0._State_3\;
                        
                    when \Quire Quire::op_OnesComplement(Quire).0._State_3\ => 
                        
                        
                        \Quire Quire::op_OnesComplement(Quire).0.binaryOperationResult.0\ := signed(SmartResize((\Quire Quire::op_OnesComplement(Quire).0.num\), 32)) < signed(SmartResize((\Quire Quire::op_OnesComplement(Quire).0.q\.\SegmentCount\), 32));
                        if (\Quire Quire::op_OnesComplement(Quire).0.binaryOperationResult.0\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Quire::op_OnesComplement(Quire).0.unaryOperationResult.0\ := not(\Quire Quire::op_OnesComplement(Quire).0.q\.\Segments\(to_integer(\Quire Quire::op_OnesComplement(Quire).0.num\)));
                            \Quire Quire::op_OnesComplement(Quire).0.q\.\Segments\(to_integer(\Quire Quire::op_OnesComplement(Quire).0.num\)) := \Quire Quire::op_OnesComplement(Quire).0.unaryOperationResult.0\;
                            
                            
                            
                            \Quire Quire::op_OnesComplement(Quire).0._State\ := \Quire Quire::op_OnesComplement(Quire).0._State_5\;
                        else 
                            \Quire Quire::op_OnesComplement(Quire).0._State\ := \Quire Quire::op_OnesComplement(Quire).0._State_4\;
                        end if;
                        
                    when \Quire Quire::op_OnesComplement(Quire).0._State_4\ => 
                        
                        
                        
                        
                        \Quire Quire::op_OnesComplement(Quire).0.return\ <= \Quire Quire::op_OnesComplement(Quire).0.q\;
                        \Quire Quire::op_OnesComplement(Quire).0._State\ := \Quire Quire::op_OnesComplement(Quire).0._State_1\;
                        
                    when \Quire Quire::op_OnesComplement(Quire).0._State_5\ => 
                        
                        \Quire Quire::op_OnesComplement(Quire).0.binaryOperationResult.1\ := SmartResize(unsigned(signed(SmartResize((\Quire Quire::op_OnesComplement(Quire).0.num\), 32)) + to_signed(1, 32)), 16);
                        \Quire Quire::op_OnesComplement(Quire).0.num\ := (\Quire Quire::op_OnesComplement(Quire).0.binaryOperationResult.1\);
                        
                        if (\Quire Quire::op_OnesComplement(Quire).0._State\ = \Quire Quire::op_OnesComplement(Quire).0._State_5\) then 
                            \Quire Quire::op_OnesComplement(Quire).0._State\ := \Quire Quire::op_OnesComplement(Quire).0._State_3\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Boolean Quire::op_Equality(Quire,Quire).0._StateMachine\: process (\Clock\) 
        Variable \Boolean Quire::op_Equality(Quire,Quire).0._State\: \Boolean Quire::op_Equality(Quire,Quire).0._States\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_0\;
        Variable \Boolean Quire::op_Equality(Quire,Quire).0.left\: \Lombiq.Arithmetics.Quire\;
        Variable \Boolean Quire::op_Equality(Quire,Quire).0.right\: \Lombiq.Arithmetics.Quire\;
        Variable \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.0\: boolean := false;
        Variable \Boolean Quire::op_Equality(Quire,Quire).0.num\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.1\: boolean := false;
        Variable \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.2\: boolean := false;
        Variable \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.3\: unsigned(15 downto 0) := to_unsigned(0, 16);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Boolean Quire::op_Equality(Quire,Quire).0._Finished\ <= false;
                \Boolean Quire::op_Equality(Quire,Quire).0.return\ <= false;
                \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_0\;
                \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.0\ := false;
                \Boolean Quire::op_Equality(Quire,Quire).0.num\ := to_unsigned(0, 16);
                \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.1\ := false;
                \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.2\ := false;
                \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.3\ := to_unsigned(0, 16);
            else 
                case \Boolean Quire::op_Equality(Quire,Quire).0._State\ is 
                    when \Boolean Quire::op_Equality(Quire,Quire).0._State_0\ => 
                        
                        
                        if (\Boolean Quire::op_Equality(Quire,Quire).0._Started\ = true) then 
                            \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_2\;
                        end if;
                        
                    when \Boolean Quire::op_Equality(Quire,Quire).0._State_1\ => 
                        
                        
                        if (\Boolean Quire::op_Equality(Quire,Quire).0._Started\ = true) then 
                            \Boolean Quire::op_Equality(Quire,Quire).0._Finished\ <= true;
                        else 
                            \Boolean Quire::op_Equality(Quire,Quire).0._Finished\ <= false;
                            \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_0\;
                        end if;
                        
                        \Boolean Quire::op_Equality(Quire,Quire).0.left.parameter.Out\ <= \Boolean Quire::op_Equality(Quire,Quire).0.left\;
                        \Boolean Quire::op_Equality(Quire,Quire).0.right.parameter.Out\ <= \Boolean Quire::op_Equality(Quire,Quire).0.right\;
                        
                    when \Boolean Quire::op_Equality(Quire,Quire).0._State_2\ => 
                        \Boolean Quire::op_Equality(Quire,Quire).0.left\ := \Boolean Quire::op_Equality(Quire,Quire).0.left.parameter.In\;
                        \Boolean Quire::op_Equality(Quire,Quire).0.right\ := \Boolean Quire::op_Equality(Quire,Quire).0.right.parameter.In\;
                        
                        
                        
                        
                        
                        \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.0\ := signed(SmartResize((\Boolean Quire::op_Equality(Quire,Quire).0.left\.\SegmentCount\), 32)) /= signed(SmartResize((\Boolean Quire::op_Equality(Quire,Quire).0.right\.\SegmentCount\), 32));

                        
                        
                        

                        if (\Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.0\) then 
                            \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_4\;
                        else 
                            
                            \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_3\;
                        end if;
                        
                    when \Boolean Quire::op_Equality(Quire,Quire).0._State_3\ => 
                        
                        
                        
                        
                        
                        
                        
                        \Boolean Quire::op_Equality(Quire,Quire).0.num\ := SmartResize(unsigned(to_signed(0, 32)), 16);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_5\;
                        
                    when \Boolean Quire::op_Equality(Quire,Quire).0._State_4\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Boolean Quire::op_Equality(Quire,Quire).0.return\ <= false;
                        \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_1\;
                        
                        if (\Boolean Quire::op_Equality(Quire,Quire).0._State\ = \Boolean Quire::op_Equality(Quire,Quire).0._State_4\) then 
                            \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_3\;
                        end if;
                        
                    when \Boolean Quire::op_Equality(Quire,Quire).0._State_5\ => 
                        
                        
                        \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.1\ := signed(SmartResize((\Boolean Quire::op_Equality(Quire,Quire).0.num\), 32)) < signed(SmartResize((\Boolean Quire::op_Equality(Quire,Quire).0.left\.\SegmentCount\), 32));
                        if (\Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.1\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.2\ := \Boolean Quire::op_Equality(Quire,Quire).0.left\.\Segments\(to_integer(\Boolean Quire::op_Equality(Quire,Quire).0.num\)) /= \Boolean Quire::op_Equality(Quire,Quire).0.right\.\Segments\(to_integer(\Boolean Quire::op_Equality(Quire,Quire).0.num\));

                            
                            
                            

                            if (\Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.2\) then 
                                \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_8\;
                            else 
                                
                                \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_7\;
                            end if;
                        else 
                            \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_6\;
                        end if;
                        
                    when \Boolean Quire::op_Equality(Quire,Quire).0._State_6\ => 
                        
                        
                        
                        
                        \Boolean Quire::op_Equality(Quire,Quire).0.return\ <= true;
                        \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_1\;
                        
                    when \Boolean Quire::op_Equality(Quire,Quire).0._State_7\ => 
                        
                        
                        
                        
                        \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.3\ := SmartResize(unsigned(signed(SmartResize((\Boolean Quire::op_Equality(Quire,Quire).0.num\), 32)) + to_signed(1, 32)), 16);
                        \Boolean Quire::op_Equality(Quire,Quire).0.num\ := (\Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.3\);
                        
                        if (\Boolean Quire::op_Equality(Quire,Quire).0._State\ = \Boolean Quire::op_Equality(Quire,Quire).0._State_7\) then 
                            \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_5\;
                        end if;
                        
                    when \Boolean Quire::op_Equality(Quire,Quire).0._State_8\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Boolean Quire::op_Equality(Quire,Quire).0.return\ <= false;
                        \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_1\;
                        
                        if (\Boolean Quire::op_Equality(Quire,Quire).0._State\ = \Boolean Quire::op_Equality(Quire,Quire).0._State_8\) then 
                            \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_7\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Quire Quire::op_RightShift(Quire,Int32).0._StateMachine\: process (\Clock\) 
        Variable \Quire Quire::op_RightShift(Quire,Int32).0._State\: \Quire Quire::op_RightShift(Quire,Int32).0._States\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_0\;
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.left\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.right\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.3\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.num\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.array\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.num2\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.4\: boolean := false;
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.flag\: boolean := false;
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.num3\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.5\: boolean := false;
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.num4\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.6\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.flag2\: boolean := false;
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.7\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.8\: boolean := false;
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.9\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.10\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.11\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.12\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.object157c924d312931f99624f9990346efe22383342001d9935b6c35c3ad8da224b8\: \Lombiq.Arithmetics.Quire\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Quire Quire::op_RightShift(Quire,Int32).0._Finished\ <= false;
                \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 64));
                \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= false;
                \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_0\;
                \Quire Quire::op_RightShift(Quire,Int32).0.right\ := to_signed(0, 32);
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.0\ := to_signed(0, 32);
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.1\ := to_signed(0, 32);
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.2\ := to_signed(0, 32);
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.3\ := to_signed(0, 32);
                \Quire Quire::op_RightShift(Quire,Int32).0.num\ := to_unsigned(0, 64);
                \Quire Quire::op_RightShift(Quire,Int32).0.array\ := (others => to_unsigned(0, 64));
                \Quire Quire::op_RightShift(Quire,Int32).0.num2\ := to_unsigned(0, 16);
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.4\ := false;
                \Quire Quire::op_RightShift(Quire,Int32).0.flag\ := false;
                \Quire Quire::op_RightShift(Quire,Int32).0.num3\ := to_unsigned(0, 16);
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.5\ := false;
                \Quire Quire::op_RightShift(Quire,Int32).0.num4\ := to_unsigned(0, 16);
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.6\ := to_unsigned(0, 16);
                \Quire Quire::op_RightShift(Quire,Int32).0.flag2\ := false;
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.7\ := to_unsigned(0, 64);
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.8\ := false;
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.9\ := to_unsigned(0, 64);
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.10\ := to_unsigned(0, 64);
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.11\ := to_unsigned(0, 16);
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.12\ := to_unsigned(0, 16);
            else 
                case \Quire Quire::op_RightShift(Quire,Int32).0._State\ is 
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_0\ => 
                        
                        
                        if (\Quire Quire::op_RightShift(Quire,Int32).0._Started\ = true) then 
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_2\;
                        end if;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_1\ => 
                        
                        
                        if (\Quire Quire::op_RightShift(Quire,Int32).0._Started\ = true) then 
                            \Quire Quire::op_RightShift(Quire,Int32).0._Finished\ <= true;
                        else 
                            \Quire Quire::op_RightShift(Quire,Int32).0._Finished\ <= false;
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_0\;
                        end if;
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.left.parameter.Out\ <= \Quire Quire::op_RightShift(Quire,Int32).0.left\;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_2\ => 
                        \Quire Quire::op_RightShift(Quire,Int32).0.left\ := \Quire Quire::op_RightShift(Quire,Int32).0.left.parameter.In\;
                        \Quire Quire::op_RightShift(Quire,Int32).0.right\ := \Quire Quire::op_RightShift(Quire,Int32).0.right.parameter.In\;
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.0\ := SmartResize(signed(SmartResize((\Quire Quire::op_RightShift(Quire,Int32).0.left\.\SegmentCount\), 32)) * to_signed(6, 32), 32);
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.1\ := shift_left(to_signed(1, 32), to_integer(unsigned(SmartResize(\Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.0\, 5))));
                        \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_3\;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_3\ => 
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.2\ := (\Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.1\) - to_signed(1, 32);
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.3\ := \Quire Quire::op_RightShift(Quire,Int32).0.right\ and (\Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.2\);
                        \Quire Quire::op_RightShift(Quire,Int32).0.right\ := \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.3\;
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.num\ := "1000000000000000000000000000000000000000000000000000000000000000";
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.array\ := (others => to_unsigned(0, 64));
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.array\ := \Quire Quire::op_RightShift(Quire,Int32).0.left\.\Segments\(0 to 7);
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.num2\ := SmartResize(unsigned(to_signed(0, 32)), 16);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_4\;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_4\ => 
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.4\ := signed(SmartResize((\Quire Quire::op_RightShift(Quire,Int32).0.num2\), 32)) < (\Quire Quire::op_RightShift(Quire,Int32).0.right\);
                        if (\Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.4\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Quire::op_RightShift(Quire,Int32).0.flag\ := false;
                            
                            
                            
                            
                            
                            
                            \Quire Quire::op_RightShift(Quire,Int32).0.num3\ := SmartResize(unsigned(to_signed(1, 32)), 16);
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_6\;
                        else 
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_5\;
                        end if;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_5\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.object157c924d312931f99624f9990346efe22383342001d9935b6c35c3ad8da224b8\.\IsNull\ := false;
                        \Quire Quire::op_RightShift(Quire,Int32).0.object157c924d312931f99624f9990346efe22383342001d9935b6c35c3ad8da224b8\.\Size\ := to_unsigned(0, 16);
                        \Quire Quire::op_RightShift(Quire,Int32).0.object157c924d312931f99624f9990346efe22383342001d9935b6c35c3ad8da224b8\.\SegmentCount\ := to_unsigned(0, 16);
                        \Quire Quire::op_RightShift(Quire,Int32).0.object157c924d312931f99624f9990346efe22383342001d9935b6c35c3ad8da224b8\.\Segments\ := (others => to_unsigned(0, 64));
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\ <= \Quire Quire::op_RightShift(Quire,Int32).0.object157c924d312931f99624f9990346efe22383342001d9935b6c35c3ad8da224b8\;
                        \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\ <= \Quire Quire::op_RightShift(Quire,Int32).0.array\;
                        \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\ <= SmartResize(unsigned(to_signed(0, 32)), 16);
                        \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= true;
                        \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_12\;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_6\ => 
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.5\ := signed(SmartResize((\Quire Quire::op_RightShift(Quire,Int32).0.num3\), 32)) <= to_signed(8, 32);
                        if (\Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.5\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.6\ := SmartResize(unsigned(to_signed(8, 32) - signed(SmartResize((\Quire Quire::op_RightShift(Quire,Int32).0.num3\), 32))), 16);
                            \Quire Quire::op_RightShift(Quire,Int32).0.num4\ := (\Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.6\);
                            
                            
                            
                            
                            
                            
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_8\;
                        else 
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_7\;
                        end if;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_7\ => 
                        
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.12\ := SmartResize(unsigned(signed(SmartResize((\Quire Quire::op_RightShift(Quire,Int32).0.num2\), 32)) + to_signed(1, 32)), 16);
                        \Quire Quire::op_RightShift(Quire,Int32).0.num2\ := (\Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.12\);
                        
                        if (\Quire Quire::op_RightShift(Quire,Int32).0._State\ = \Quire Quire::op_RightShift(Quire,Int32).0._State_7\) then 
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_4\;
                        end if;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_8\ => 
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.7\ := \Quire Quire::op_RightShift(Quire,Int32).0.array\(to_integer(\Quire Quire::op_RightShift(Quire,Int32).0.num4\)) and to_unsigned(1, 64);
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.8\ := (\Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.7\) = to_unsigned(1, 64);
                        \Quire Quire::op_RightShift(Quire,Int32).0.flag2\ := \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.8\;
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_9\;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_9\ => 
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.9\ := SmartResize(shift_right(\Quire Quire::op_RightShift(Quire,Int32).0.array\(to_integer(\Quire Quire::op_RightShift(Quire,Int32).0.num4\)), to_integer(unsigned(SmartResize(to_signed(1, 32), 6) and "111111"))), 64);
                        \Quire Quire::op_RightShift(Quire,Int32).0.array\(to_integer(\Quire Quire::op_RightShift(Quire,Int32).0.num4\)) := \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.9\;
                        
                        
                        
                        
                        

                        
                        
                        

                        if (\Quire Quire::op_RightShift(Quire,Int32).0.flag\) then 
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_11\;
                        else 
                            
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_10\;
                        end if;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_10\ => 
                        
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.flag\ := \Quire Quire::op_RightShift(Quire,Int32).0.flag2\;
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.11\ := SmartResize(unsigned(signed(SmartResize((\Quire Quire::op_RightShift(Quire,Int32).0.num3\), 32)) + to_signed(1, 32)), 16);
                        \Quire Quire::op_RightShift(Quire,Int32).0.num3\ := (\Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.11\);
                        
                        if (\Quire Quire::op_RightShift(Quire,Int32).0._State\ = \Quire Quire::op_RightShift(Quire,Int32).0._State_10\) then 
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_6\;
                        end if;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_11\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.10\ := \Quire Quire::op_RightShift(Quire,Int32).0.array\(to_integer(\Quire Quire::op_RightShift(Quire,Int32).0.num4\)) or \Quire Quire::op_RightShift(Quire,Int32).0.num\;
                        \Quire Quire::op_RightShift(Quire,Int32).0.array\(to_integer(\Quire Quire::op_RightShift(Quire,Int32).0.num4\)) := \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.10\;
                        
                        if (\Quire Quire::op_RightShift(Quire,Int32).0._State\ = \Quire Quire::op_RightShift(Quire,Int32).0._State_11\) then 
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_10\;
                        end if;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_12\ => 
                        
                        if (\Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ = \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\) then 
                            \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= false;
                            \Quire Quire::op_RightShift(Quire,Int32).0.object157c924d312931f99624f9990346efe22383342001d9935b6c35c3ad8da224b8\ := \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\;
                            \Quire Quire::op_RightShift(Quire,Int32).0.array\ := \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\;
                            
                            
                            
                            \Quire Quire::op_RightShift(Quire,Int32).0.return\ <= \Quire Quire::op_RightShift(Quire,Int32).0.object157c924d312931f99624f9990346efe22383342001d9935b6c35c3ad8da224b8\;
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_1\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Quire Quire::op_LeftShift(Quire,Int32).0._StateMachine\: process (\Clock\) 
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0._State\: \Quire Quire::op_LeftShift(Quire,Int32).0._States\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_0\;
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.left\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.right\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.num\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.array\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.num2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.num3\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.1\: boolean := false;
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.flag\: boolean := false;
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.num4\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.2\: boolean := false;
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.flag2\: boolean := false;
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.3\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.4\: boolean := false;
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.5\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.6\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.7\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.8\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.objectc996901721b3380940539d5e2ccc153d36bc5159fbc7657e5cc431d1b5e93c1f\: \Lombiq.Arithmetics.Quire\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Quire Quire::op_LeftShift(Quire,Int32).0._Finished\ <= false;
                \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 64));
                \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= false;
                \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_0\;
                \Quire Quire::op_LeftShift(Quire,Int32).0.right\ := to_signed(0, 32);
                \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.0\ := to_signed(0, 32);
                \Quire Quire::op_LeftShift(Quire,Int32).0.num\ := to_unsigned(0, 64);
                \Quire Quire::op_LeftShift(Quire,Int32).0.array\ := (others => to_unsigned(0, 64));
                \Quire Quire::op_LeftShift(Quire,Int32).0.num2\ := to_unsigned(0, 32);
                \Quire Quire::op_LeftShift(Quire,Int32).0.num3\ := to_unsigned(0, 16);
                \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.1\ := false;
                \Quire Quire::op_LeftShift(Quire,Int32).0.flag\ := false;
                \Quire Quire::op_LeftShift(Quire,Int32).0.num4\ := to_unsigned(0, 16);
                \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.2\ := false;
                \Quire Quire::op_LeftShift(Quire,Int32).0.flag2\ := false;
                \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.3\ := to_unsigned(0, 64);
                \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.4\ := false;
                \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.5\ := to_unsigned(0, 64);
                \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.6\ := to_unsigned(0, 64);
                \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.7\ := to_unsigned(0, 16);
                \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.8\ := to_unsigned(0, 16);
            else 
                case \Quire Quire::op_LeftShift(Quire,Int32).0._State\ is 
                    when \Quire Quire::op_LeftShift(Quire,Int32).0._State_0\ => 
                        
                        
                        if (\Quire Quire::op_LeftShift(Quire,Int32).0._Started\ = true) then 
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_2\;
                        end if;
                        
                    when \Quire Quire::op_LeftShift(Quire,Int32).0._State_1\ => 
                        
                        
                        if (\Quire Quire::op_LeftShift(Quire,Int32).0._Started\ = true) then 
                            \Quire Quire::op_LeftShift(Quire,Int32).0._Finished\ <= true;
                        else 
                            \Quire Quire::op_LeftShift(Quire,Int32).0._Finished\ <= false;
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_0\;
                        end if;
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.left.parameter.Out\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.left\;
                        
                    when \Quire Quire::op_LeftShift(Quire,Int32).0._State_2\ => 
                        \Quire Quire::op_LeftShift(Quire,Int32).0.left\ := \Quire Quire::op_LeftShift(Quire,Int32).0.left.parameter.In\;
                        \Quire Quire::op_LeftShift(Quire,Int32).0.right\ := \Quire Quire::op_LeftShift(Quire,Int32).0.right.parameter.In\;
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.0\ := \Quire Quire::op_LeftShift(Quire,Int32).0.right\ and to_signed(65535, 32);
                        \Quire Quire::op_LeftShift(Quire,Int32).0.right\ := \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.0\;
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.num\ := "1000000000000000000000000000000000000000000000000000000000000000";
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.array\ := (others => to_unsigned(0, 64));
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.array\ := \Quire Quire::op_LeftShift(Quire,Int32).0.left\.\Segments\(0 to 7);
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.num2\ := to_unsigned(1, 32);
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.num3\ := SmartResize(unsigned(to_signed(0, 32)), 16);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_3\;
                        
                    when \Quire Quire::op_LeftShift(Quire,Int32).0._State_3\ => 
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.1\ := signed(SmartResize((\Quire Quire::op_LeftShift(Quire,Int32).0.num3\), 32)) < (\Quire Quire::op_LeftShift(Quire,Int32).0.right\);
                        if (\Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.1\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Quire::op_LeftShift(Quire,Int32).0.flag\ := false;
                            
                            
                            
                            
                            
                            
                            \Quire Quire::op_LeftShift(Quire,Int32).0.num4\ := SmartResize(unsigned(to_signed(0, 32)), 16);
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_5\;
                        else 
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_4\;
                        end if;
                        
                    when \Quire Quire::op_LeftShift(Quire,Int32).0._State_4\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.objectc996901721b3380940539d5e2ccc153d36bc5159fbc7657e5cc431d1b5e93c1f\.\IsNull\ := false;
                        \Quire Quire::op_LeftShift(Quire,Int32).0.objectc996901721b3380940539d5e2ccc153d36bc5159fbc7657e5cc431d1b5e93c1f\.\Size\ := to_unsigned(0, 16);
                        \Quire Quire::op_LeftShift(Quire,Int32).0.objectc996901721b3380940539d5e2ccc153d36bc5159fbc7657e5cc431d1b5e93c1f\.\SegmentCount\ := to_unsigned(0, 16);
                        \Quire Quire::op_LeftShift(Quire,Int32).0.objectc996901721b3380940539d5e2ccc153d36bc5159fbc7657e5cc431d1b5e93c1f\.\Segments\ := (others => to_unsigned(0, 64));
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.objectc996901721b3380940539d5e2ccc153d36bc5159fbc7657e5cc431d1b5e93c1f\;
                        \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.array\;
                        \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\ <= SmartResize(unsigned(to_signed(0, 32)), 16);
                        \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= true;
                        \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_10\;
                        
                    when \Quire Quire::op_LeftShift(Quire,Int32).0._State_5\ => 
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.2\ := signed(SmartResize((\Quire Quire::op_LeftShift(Quire,Int32).0.num4\), 32)) < to_signed(8, 32);
                        if (\Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.2\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.3\ := \Quire Quire::op_LeftShift(Quire,Int32).0.array\(to_integer(\Quire Quire::op_LeftShift(Quire,Int32).0.num4\)) and \Quire Quire::op_LeftShift(Quire,Int32).0.num\;
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_7\;
                        else 
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_6\;
                        end if;
                        
                    when \Quire Quire::op_LeftShift(Quire,Int32).0._State_6\ => 
                        
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.8\ := SmartResize(unsigned(signed(SmartResize((\Quire Quire::op_LeftShift(Quire,Int32).0.num3\), 32)) + to_signed(1, 32)), 16);
                        \Quire Quire::op_LeftShift(Quire,Int32).0.num3\ := (\Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.8\);
                        
                        if (\Quire Quire::op_LeftShift(Quire,Int32).0._State\ = \Quire Quire::op_LeftShift(Quire,Int32).0._State_6\) then 
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_3\;
                        end if;
                        
                    when \Quire Quire::op_LeftShift(Quire,Int32).0._State_7\ => 
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.4\ := (\Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.3\) = \Quire Quire::op_LeftShift(Quire,Int32).0.num\;
                        \Quire Quire::op_LeftShift(Quire,Int32).0.flag2\ := \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.4\;
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.5\ := SmartResize(shift_left(\Quire Quire::op_LeftShift(Quire,Int32).0.array\(to_integer(\Quire Quire::op_LeftShift(Quire,Int32).0.num4\)), to_integer(unsigned(SmartResize(to_signed(1, 32), 6)))), 64);
                        \Quire Quire::op_LeftShift(Quire,Int32).0.array\(to_integer(\Quire Quire::op_LeftShift(Quire,Int32).0.num4\)) := \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.5\;
                        
                        
                        
                        
                        

                        
                        
                        

                        if (\Quire Quire::op_LeftShift(Quire,Int32).0.flag\) then 
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_9\;
                        else 
                            
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_8\;
                        end if;
                        
                    when \Quire Quire::op_LeftShift(Quire,Int32).0._State_8\ => 
                        
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.flag\ := \Quire Quire::op_LeftShift(Quire,Int32).0.flag2\;
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.7\ := SmartResize(unsigned(signed(SmartResize((\Quire Quire::op_LeftShift(Quire,Int32).0.num4\), 32)) + to_signed(1, 32)), 16);
                        \Quire Quire::op_LeftShift(Quire,Int32).0.num4\ := (\Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.7\);
                        
                        if (\Quire Quire::op_LeftShift(Quire,Int32).0._State\ = \Quire Quire::op_LeftShift(Quire,Int32).0._State_8\) then 
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_5\;
                        end if;
                        
                    when \Quire Quire::op_LeftShift(Quire,Int32).0._State_9\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.6\ := \Quire Quire::op_LeftShift(Quire,Int32).0.array\(to_integer(\Quire Quire::op_LeftShift(Quire,Int32).0.num4\)) or SmartResize((\Quire Quire::op_LeftShift(Quire,Int32).0.num2\), 64);
                        \Quire Quire::op_LeftShift(Quire,Int32).0.array\(to_integer(\Quire Quire::op_LeftShift(Quire,Int32).0.num4\)) := (\Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.6\);
                        
                        if (\Quire Quire::op_LeftShift(Quire,Int32).0._State\ = \Quire Quire::op_LeftShift(Quire,Int32).0._State_9\) then 
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_8\;
                        end if;
                        
                    when \Quire Quire::op_LeftShift(Quire,Int32).0._State_10\ => 
                        
                        if (\Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ = \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\) then 
                            \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= false;
                            \Quire Quire::op_LeftShift(Quire,Int32).0.objectc996901721b3380940539d5e2ccc153d36bc5159fbc7657e5cc431d1b5e93c1f\ := \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\;
                            \Quire Quire::op_LeftShift(Quire,Int32).0.array\ := \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\;
                            
                            
                            
                            \Quire Quire::op_LeftShift(Quire,Int32).0.return\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.objectc996901721b3380940539d5e2ccc153d36bc5159fbc7657e5cc431d1b5e93c1f\;
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_1\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \UInt64 Quire::op_Explicit(Quire).0._StateMachine\: process (\Clock\) 
        Variable \UInt64 Quire::op_Explicit(Quire).0._State\: \UInt64 Quire::op_Explicit(Quire).0._States\ := \UInt64 Quire::op_Explicit(Quire).0._State_0\;
        Variable \UInt64 Quire::op_Explicit(Quire).0.x\: \Lombiq.Arithmetics.Quire\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \UInt64 Quire::op_Explicit(Quire).0._Finished\ <= false;
                \UInt64 Quire::op_Explicit(Quire).0.return\ <= to_unsigned(0, 64);
                \UInt64 Quire::op_Explicit(Quire).0._State\ := \UInt64 Quire::op_Explicit(Quire).0._State_0\;
            else 
                case \UInt64 Quire::op_Explicit(Quire).0._State\ is 
                    when \UInt64 Quire::op_Explicit(Quire).0._State_0\ => 
                        
                        
                        if (\UInt64 Quire::op_Explicit(Quire).0._Started\ = true) then 
                            \UInt64 Quire::op_Explicit(Quire).0._State\ := \UInt64 Quire::op_Explicit(Quire).0._State_2\;
                        end if;
                        
                    when \UInt64 Quire::op_Explicit(Quire).0._State_1\ => 
                        
                        
                        if (\UInt64 Quire::op_Explicit(Quire).0._Started\ = true) then 
                            \UInt64 Quire::op_Explicit(Quire).0._Finished\ <= true;
                        else 
                            \UInt64 Quire::op_Explicit(Quire).0._Finished\ <= false;
                            \UInt64 Quire::op_Explicit(Quire).0._State\ := \UInt64 Quire::op_Explicit(Quire).0._State_0\;
                        end if;
                        
                        \UInt64 Quire::op_Explicit(Quire).0.x.parameter.Out\ <= \UInt64 Quire::op_Explicit(Quire).0.x\;
                        
                    when \UInt64 Quire::op_Explicit(Quire).0._State_2\ => 
                        \UInt64 Quire::op_Explicit(Quire).0.x\ := \UInt64 Quire::op_Explicit(Quire).0.x.parameter.In\;
                        
                        
                        
                        \UInt64 Quire::op_Explicit(Quire).0.return\ <= \UInt64 Quire::op_Explicit(Quire).0.x\.\Segments\(to_integer(to_signed(0, 32)));
                        \UInt64 Quire::op_Explicit(Quire).0._State\ := \UInt64 Quire::op_Explicit(Quire).0._State_1\;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \UInt32 Quire::op_Explicit(Quire).0._StateMachine\: process (\Clock\) 
        Variable \UInt32 Quire::op_Explicit(Quire).0._State\: \UInt32 Quire::op_Explicit(Quire).0._States\ := \UInt32 Quire::op_Explicit(Quire).0._State_0\;
        Variable \UInt32 Quire::op_Explicit(Quire).0.x\: \Lombiq.Arithmetics.Quire\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \UInt32 Quire::op_Explicit(Quire).0._Finished\ <= false;
                \UInt32 Quire::op_Explicit(Quire).0.return\ <= to_unsigned(0, 32);
                \UInt32 Quire::op_Explicit(Quire).0._State\ := \UInt32 Quire::op_Explicit(Quire).0._State_0\;
            else 
                case \UInt32 Quire::op_Explicit(Quire).0._State\ is 
                    when \UInt32 Quire::op_Explicit(Quire).0._State_0\ => 
                        
                        
                        if (\UInt32 Quire::op_Explicit(Quire).0._Started\ = true) then 
                            \UInt32 Quire::op_Explicit(Quire).0._State\ := \UInt32 Quire::op_Explicit(Quire).0._State_2\;
                        end if;
                        
                    when \UInt32 Quire::op_Explicit(Quire).0._State_1\ => 
                        
                        
                        if (\UInt32 Quire::op_Explicit(Quire).0._Started\ = true) then 
                            \UInt32 Quire::op_Explicit(Quire).0._Finished\ <= true;
                        else 
                            \UInt32 Quire::op_Explicit(Quire).0._Finished\ <= false;
                            \UInt32 Quire::op_Explicit(Quire).0._State\ := \UInt32 Quire::op_Explicit(Quire).0._State_0\;
                        end if;
                        
                        \UInt32 Quire::op_Explicit(Quire).0.x.parameter.Out\ <= \UInt32 Quire::op_Explicit(Quire).0.x\;
                        
                    when \UInt32 Quire::op_Explicit(Quire).0._State_2\ => 
                        \UInt32 Quire::op_Explicit(Quire).0.x\ := \UInt32 Quire::op_Explicit(Quire).0.x.parameter.In\;
                        
                        
                        
                        \UInt32 Quire::op_Explicit(Quire).0.return\ <= SmartResize(\UInt32 Quire::op_Explicit(Quire).0.x\.\Segments\(to_integer(to_signed(0, 32))), 32);
                        \UInt32 Quire::op_Explicit(Quire).0._State\ := \UInt32 Quire::op_Explicit(Quire).0._State_1\;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Finished\ <= \FinishedInternal\;
    \Hast::ExternalInvocationProxy()\: process (\Clock\) 
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \FinishedInternal\ <= false;
                \Hast::ExternalInvocationProxy().Posit32FusedCalculator::CalculateFusedSum(SimpleMemory)._Started.0\ <= false;
            else 
                if (\Started\ = true and \FinishedInternal\ = false) then 
                    
                    case \MemberId\ is 
                        when 0 => 
                            if (\Hast::ExternalInvocationProxy().Posit32FusedCalculator::CalculateFusedSum(SimpleMemory)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().Posit32FusedCalculator::CalculateFusedSum(SimpleMemory)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().Posit32FusedCalculator::CalculateFusedSum(SimpleMemory)._Started.0\ = \Hast::ExternalInvocationProxy().Posit32FusedCalculator::CalculateFusedSum(SimpleMemory)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().Posit32FusedCalculator::CalculateFusedSum(SimpleMemory)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when others => 
                            null;
                    end case;
                else 
                    
                    if (\Started\ = false and \FinishedInternal\ = true) then 
                        \FinishedInternal\ <= false;
                    end if;
                end if;
            end if;
        end if;
    end process;
    


    
    
    \Posit32::.ctor(Int32).0._Started\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Started.0\;
    \Posit32::.ctor(Int32).0.this.parameter.In\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).this.parameter.Out.0\;
    \Posit32::.ctor(Int32).0.value.parameter.In\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).value.parameter.Out.0\;
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Finished.0\ <= \Posit32::.ctor(Int32).0._Finished\;
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).this.parameter.In.0\ <= \Posit32::.ctor(Int32).0.this.parameter.Out\;
    


    
    \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForStarted;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\ <= false;
                \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\ <= false;
            else 

                
                case \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Started.0\) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.runningIndex.0\ := 0;
                            \Quire Posit32::op_Explicit(Posit32).0._Started\ <= true;
                            \Quire Posit32::op_Explicit(Posit32).0.x.parameter.In\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32).x.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire Posit32::op_Explicit(Posit32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\ <= true;
                                    \Quire Posit32::op_Explicit(Posit32).0._Started\ <= false;
                                    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32).return.0\ <= \Quire Posit32::op_Explicit(Posit32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Started.0\) then 
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ := 0;
                            \Quire Posit32::op_Explicit(Posit32).0._Started\ <= true;
                            \Quire Posit32::op_Explicit(Posit32).0.x.parameter.In\ <= \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32).x.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire Posit32::op_Explicit(Posit32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := AfterFinished;
                                    \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\ <= true;
                                    \Quire Posit32::op_Explicit(Posit32).0._Started\ <= false;
                                    \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32).return.0\ <= \Quire Posit32::op_Explicit(Posit32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForStarted;
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    


    
    
    \Posit32::.ctor(UInt32,Boolean).0._Started\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean)._Started.0\;
    \Posit32::.ctor(UInt32,Boolean).0.this.parameter.In\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).this.parameter.Out.0\;
    \Posit32::.ctor(UInt32,Boolean).0.bits.parameter.In\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).bits.parameter.Out.0\;
    \Posit32::.ctor(UInt32,Boolean).0.fromBitMask.parameter.In\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).fromBitMask.parameter.Out.0\;
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean)._Finished.0\ <= \Posit32::.ctor(UInt32,Boolean).0._Finished\;
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).this.parameter.In.0\ <= \Posit32::.ctor(UInt32,Boolean).0.this.parameter.Out\;
    


    
    
    \Posit32::FusedSum(Posit32[],Quire).0._Started\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire)._Started.0\;
    \Posit32::FusedSum(Posit32[],Quire).0.posits.parameter.In\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).posits.parameter.Out.0\;
    \Posit32::FusedSum(Posit32[],Quire).0.startingValue.parameter.In\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).startingValue.parameter.Out.0\;
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire)._Finished.0\ <= \Posit32::FusedSum(Posit32[],Quire).0._Finished\;
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).return.0\ <= \Posit32::FusedSum(Posit32[],Quire).0.return\;
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).posits.parameter.In.0\ <= \Posit32::FusedSum(Posit32[],Quire).0.posits.parameter.Out\;
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).startingValue.parameter.In.0\ <= \Posit32::FusedSum(Posit32[],Quire).0.startingValue.parameter.Out\;
    


    
    
    \Posit32::.ctor(Quire).0._Started\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire)._Started.0\;
    \Posit32::.ctor(Quire).0.this.parameter.In\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).this.parameter.Out.0\;
    \Posit32::.ctor(Quire).0.q.parameter.In\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).q.parameter.Out.0\;
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire)._Finished.0\ <= \Posit32::.ctor(Quire).0._Finished\;
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).this.parameter.In.0\ <= \Posit32::.ctor(Quire).0.this.parameter.Out\;
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).q.parameter.In.0\ <= \Posit32::.ctor(Quire).0.q.parameter.Out\;
    


    
    
    \Quire Quire::op_RightShift(Quire,Int32).0._Started\ <= \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\;
    \Quire Quire::op_RightShift(Quire,Int32).0.left.parameter.In\ <= \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.Out.0\;
    \Quire Quire::op_RightShift(Quire,Int32).0.right.parameter.In\ <= \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).right.parameter.Out.0\;
    \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Finished.0\ <= \Quire Quire::op_RightShift(Quire,Int32).0._Finished\;
    \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).return.0\ <= \Quire Quire::op_RightShift(Quire,Int32).0.return\;
    \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.In.0\ <= \Quire Quire::op_RightShift(Quire,Int32).0.left.parameter.Out\;
    


    
    
    \UInt64 Quire::op_Explicit(Quire).0._Started\ <= \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\;
    \UInt64 Quire::op_Explicit(Quire).0.x.parameter.In\ <= \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).x.parameter.Out.0\;
    \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Finished.0\ <= \UInt64 Quire::op_Explicit(Quire).0._Finished\;
    \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).return.0\ <= \UInt64 Quire::op_Explicit(Quire).0.return\;
    \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).x.parameter.In.0\ <= \UInt64 Quire::op_Explicit(Quire).0.x.parameter.Out\;
    


    
    
    \Quire Quire::op_OnesComplement(Quire).0._Started\ <= \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire)._Started.0\;
    \Quire Quire::op_OnesComplement(Quire).0.q.parameter.In\ <= \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire).q.parameter.Out.0\;
    \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire)._Finished.0\ <= \Quire Quire::op_OnesComplement(Quire).0._Finished\;
    \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire).return.0\ <= \Quire Quire::op_OnesComplement(Quire).0.return\;
    \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire).q.parameter.In.0\ <= \Quire Quire::op_OnesComplement(Quire).0.q.parameter.Out\;
    


    
    
    \Quire Quire::op_Addition(Quire,UInt32).0._Started\ <= \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32)._Started.0\;
    \Quire Quire::op_Addition(Quire,UInt32).0.left.parameter.In\ <= \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).left.parameter.Out.0\;
    \Quire Quire::op_Addition(Quire,UInt32).0.right.parameter.In\ <= \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).right.parameter.Out.0\;
    \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32)._Finished.0\ <= \Quire Quire::op_Addition(Quire,UInt32).0._Finished\;
    \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).return.0\ <= \Quire Quire::op_Addition(Quire,UInt32).0.return\;
    \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).left.parameter.In.0\ <= \Quire Quire::op_Addition(Quire,UInt32).0.left.parameter.Out\;
    


    
    \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::.ctor(Quire).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::.ctor(Quire).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Quire Posit32::op_Explicit(Posit32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::.ctor(Quire).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::.ctor(Quire).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForStarted;
                \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= false;
                \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= false;
                \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= false;
            else 

                
                case \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::.ctor(Quire).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\) then 
                            \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::.ctor(Quire).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::.ctor(Quire).0.runningIndex.0\ := 0;
                            \Quire Quire::op_LeftShift(Quire,Int32).0._Started\ <= true;
                            \Quire Quire::op_LeftShift(Quire,Int32).0.left.parameter.In\ <= \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.Out.0\;
                            \Quire Quire::op_LeftShift(Quire,Int32).0.right.parameter.In\ <= \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::.ctor(Quire).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire Quire::op_LeftShift(Quire,Int32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::.ctor(Quire).0.runningState.0\ := AfterFinished;
                                    \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= true;
                                    \Quire Quire::op_LeftShift(Quire,Int32).0._Started\ <= false;
                                    \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).return.0\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.return\;
                                    \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.In.0\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.left.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::.ctor(Quire).0.runningState.0\ := WaitingForStarted;
                            \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\) then 
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ := 0;
                            \Quire Quire::op_LeftShift(Quire,Int32).0._Started\ <= true;
                            \Quire Quire::op_LeftShift(Quire,Int32).0.left.parameter.In\ <= \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.Out.0\;
                            \Quire Quire::op_LeftShift(Quire,Int32).0.right.parameter.In\ <= \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire Quire::op_LeftShift(Quire,Int32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := AfterFinished;
                                    \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= true;
                                    \Quire Quire::op_LeftShift(Quire,Int32).0._Started\ <= false;
                                    \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).return.0\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.return\;
                                    \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.In.0\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.left.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForStarted;
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\) then 
                            \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ := 0;
                            \Quire Quire::op_LeftShift(Quire,Int32).0._Started\ <= true;
                            \Quire Quire::op_LeftShift(Quire,Int32).0.left.parameter.In\ <= \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.Out.0\;
                            \Quire Quire::op_LeftShift(Quire,Int32).0.right.parameter.In\ <= \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire Quire::op_LeftShift(Quire,Int32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := AfterFinished;
                                    \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= true;
                                    \Quire Quire::op_LeftShift(Quire,Int32).0._Started\ <= false;
                                    \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).return.0\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.return\;
                                    \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.In.0\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.left.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForStarted;
                            \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    


    
    
    \UInt32 Quire::op_Explicit(Quire).0._Started\ <= \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire)._Started.0\;
    \UInt32 Quire::op_Explicit(Quire).0.x.parameter.In\ <= \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire).x.parameter.Out.0\;
    \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire)._Finished.0\ <= \UInt32 Quire::op_Explicit(Quire).0._Finished\;
    \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire).return.0\ <= \UInt32 Quire::op_Explicit(Quire).0.return\;
    \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire).x.parameter.In.0\ <= \UInt32 Quire::op_Explicit(Quire).0.x.parameter.Out\;
    


    
    
    \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._Started\ <= \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32)._Started.0\;
    \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.signBit.parameter.In\ <= \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).signBit.parameter.Out.0\;
    \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.regimeKValue.parameter.In\ <= \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).regimeKValue.parameter.Out.0\;
    \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits.parameter.In\ <= \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).exponentBits.parameter.Out.0\;
    \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits.parameter.In\ <= \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).fractionBits.parameter.Out.0\;
    \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32)._Finished.0\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._Finished\;
    \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).return.0\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return\;
    


    
    
    \Posit32::.ctor(UInt32).0._Started\ <= \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32)._Started.0\;
    \Posit32::.ctor(UInt32).0.this.parameter.In\ <= \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32).this.parameter.Out.0\;
    \Posit32::.ctor(UInt32).0.value.parameter.In\ <= \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32).value.parameter.Out.0\;
    \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32)._Finished.0\ <= \Posit32::.ctor(UInt32).0._Finished\;
    \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32).this.parameter.In.0\ <= \Posit32::.ctor(UInt32).0.this.parameter.Out\;
    


    
    \Hast::InternalInvocationProxy().Posit32::GetMostSignificantOnePosition(UInt32)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Posit32::GetMostSignificantOnePosition(UInt32).Posit32::EncodeRegimeBits(Int32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Posit32::GetMostSignificantOnePosition(UInt32).Posit32::EncodeRegimeBits(Int32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Posit32::GetMostSignificantOnePosition(UInt32).Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Posit32::GetMostSignificantOnePosition(UInt32).Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Hast::InternalInvocationProxy().Posit32::GetMostSignificantOnePosition(UInt32).Posit32::EncodeRegimeBits(Int32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Posit32::GetMostSignificantOnePosition(UInt32).Posit32::EncodeRegimeBits(Int32).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Posit32::GetMostSignificantOnePosition(UInt32).Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Posit32::GetMostSignificantOnePosition(UInt32).Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.runningState.0\ := WaitingForStarted;
                \Posit32::EncodeRegimeBits(Int32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Finished.0\ <= false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Finished.0\ <= false;
            else 

                
                case \Hast::InternalInvocationProxy().Posit32::GetMostSignificantOnePosition(UInt32).Posit32::EncodeRegimeBits(Int32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Posit32::EncodeRegimeBits(Int32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Started.0\) then 
                            \Posit32::EncodeRegimeBits(Int32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Posit32::GetMostSignificantOnePosition(UInt32).Posit32::EncodeRegimeBits(Int32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Posit32::GetMostSignificantOnePosition(UInt32).Posit32::EncodeRegimeBits(Int32).0.runningIndex.0\ := 0;
                            \Posit32::GetMostSignificantOnePosition(UInt32).0._Started\ <= true;
                            \Posit32::GetMostSignificantOnePosition(UInt32).0.bits.parameter.In\ <= \Posit32::EncodeRegimeBits(Int32).0.Posit32::GetMostSignificantOnePosition(UInt32).bits.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Posit32::GetMostSignificantOnePosition(UInt32).Posit32::EncodeRegimeBits(Int32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Posit32::GetMostSignificantOnePosition(UInt32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Posit32::GetMostSignificantOnePosition(UInt32).Posit32::EncodeRegimeBits(Int32).0.runningState.0\ := AfterFinished;
                                    \Posit32::EncodeRegimeBits(Int32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Finished.0\ <= true;
                                    \Posit32::GetMostSignificantOnePosition(UInt32).0._Started\ <= false;
                                    \Posit32::EncodeRegimeBits(Int32).0.Posit32::GetMostSignificantOnePosition(UInt32).return.0\ <= \Posit32::GetMostSignificantOnePosition(UInt32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Posit32::EncodeRegimeBits(Int32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Posit32::GetMostSignificantOnePosition(UInt32).Posit32::EncodeRegimeBits(Int32).0.runningState.0\ := WaitingForStarted;
                            \Posit32::EncodeRegimeBits(Int32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Posit32::GetMostSignificantOnePosition(UInt32).Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Started.0\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Posit32::GetMostSignificantOnePosition(UInt32).Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Posit32::GetMostSignificantOnePosition(UInt32).Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.runningIndex.0\ := 0;
                            \Posit32::GetMostSignificantOnePosition(UInt32).0._Started\ <= true;
                            \Posit32::GetMostSignificantOnePosition(UInt32).0.bits.parameter.In\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetMostSignificantOnePosition(UInt32).bits.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Posit32::GetMostSignificantOnePosition(UInt32).Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Posit32::GetMostSignificantOnePosition(UInt32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Posit32::GetMostSignificantOnePosition(UInt32).Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.runningState.0\ := AfterFinished;
                                    \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Finished.0\ <= true;
                                    \Posit32::GetMostSignificantOnePosition(UInt32).0._Started\ <= false;
                                    \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetMostSignificantOnePosition(UInt32).return.0\ <= \Posit32::GetMostSignificantOnePosition(UInt32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Posit32::GetMostSignificantOnePosition(UInt32).Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.runningState.0\ := WaitingForStarted;
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetMostSignificantOnePosition(UInt32)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    


    
    
    \Posit32::EncodeRegimeBits(Int32).0._Started\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::EncodeRegimeBits(Int32)._Started.0\;
    \Posit32::EncodeRegimeBits(Int32).0.regimeKValue.parameter.In\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::EncodeRegimeBits(Int32).regimeKValue.parameter.Out.0\;
    \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::EncodeRegimeBits(Int32)._Finished.0\ <= \Posit32::EncodeRegimeBits(Int32).0._Finished\;
    \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::EncodeRegimeBits(Int32).return.0\ <= \Posit32::EncodeRegimeBits(Int32).0.return\;
    


    
    \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::GetRegimeKValue().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::GetRegimeKValue().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::ExponentSize().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::ExponentSize().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::FractionSize().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::FractionSize().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::GetRegimeKValue().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::GetRegimeKValue().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::ExponentSize().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::ExponentSize().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::FractionSize().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::FractionSize().0.runningState.0\ := WaitingForStarted;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\ <= false;
                \Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\ <= false;
                \Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\ <= false;
                \Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\ <= false;
            else 

                
                case \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.runningIndex.0\ := 0;
                            \Posit32::LengthOfRunOfBits(UInt32,Byte).0._Started\ <= true;
                            \Posit32::LengthOfRunOfBits(UInt32,Byte).0.bits.parameter.In\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte).bits.parameter.Out.0\;
                            \Posit32::LengthOfRunOfBits(UInt32,Byte).0.startingPosition.parameter.In\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte).startingPosition.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Posit32::LengthOfRunOfBits(UInt32,Byte).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.runningState.0\ := AfterFinished;
                                    \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\ <= true;
                                    \Posit32::LengthOfRunOfBits(UInt32,Byte).0._Started\ <= false;
                                    \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte).return.0\ <= \Posit32::LengthOfRunOfBits(UInt32,Byte).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.runningState.0\ := WaitingForStarted;
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::GetRegimeKValue().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\) then 
                            \Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::GetRegimeKValue().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::GetRegimeKValue().0.runningIndex.0\ := 0;
                            \Posit32::LengthOfRunOfBits(UInt32,Byte).0._Started\ <= true;
                            \Posit32::LengthOfRunOfBits(UInt32,Byte).0.bits.parameter.In\ <= \Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte).bits.parameter.Out.0\;
                            \Posit32::LengthOfRunOfBits(UInt32,Byte).0.startingPosition.parameter.In\ <= \Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte).startingPosition.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::GetRegimeKValue().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Posit32::LengthOfRunOfBits(UInt32,Byte).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::GetRegimeKValue().0.runningState.0\ := AfterFinished;
                                    \Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\ <= true;
                                    \Posit32::LengthOfRunOfBits(UInt32,Byte).0._Started\ <= false;
                                    \Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte).return.0\ <= \Posit32::LengthOfRunOfBits(UInt32,Byte).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::GetRegimeKValue().0.runningState.0\ := WaitingForStarted;
                            \Posit32::GetRegimeKValue().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::ExponentSize().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\) then 
                            \Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::ExponentSize().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::ExponentSize().0.runningIndex.0\ := 0;
                            \Posit32::LengthOfRunOfBits(UInt32,Byte).0._Started\ <= true;
                            \Posit32::LengthOfRunOfBits(UInt32,Byte).0.bits.parameter.In\ <= \Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte).bits.parameter.Out.0\;
                            \Posit32::LengthOfRunOfBits(UInt32,Byte).0.startingPosition.parameter.In\ <= \Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte).startingPosition.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::ExponentSize().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Posit32::LengthOfRunOfBits(UInt32,Byte).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::ExponentSize().0.runningState.0\ := AfterFinished;
                                    \Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\ <= true;
                                    \Posit32::LengthOfRunOfBits(UInt32,Byte).0._Started\ <= false;
                                    \Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte).return.0\ <= \Posit32::LengthOfRunOfBits(UInt32,Byte).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::ExponentSize().0.runningState.0\ := WaitingForStarted;
                            \Posit32::ExponentSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::FractionSize().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\) then 
                            \Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::FractionSize().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::FractionSize().0.runningIndex.0\ := 0;
                            \Posit32::LengthOfRunOfBits(UInt32,Byte).0._Started\ <= true;
                            \Posit32::LengthOfRunOfBits(UInt32,Byte).0.bits.parameter.In\ <= \Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte).bits.parameter.Out.0\;
                            \Posit32::LengthOfRunOfBits(UInt32,Byte).0.startingPosition.parameter.In\ <= \Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte).startingPosition.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::FractionSize().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Posit32::LengthOfRunOfBits(UInt32,Byte).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::FractionSize().0.runningState.0\ := AfterFinished;
                                    \Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\ <= true;
                                    \Posit32::LengthOfRunOfBits(UInt32,Byte).0._Started\ <= false;
                                    \Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte).return.0\ <= \Posit32::LengthOfRunOfBits(UInt32,Byte).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Posit32::LengthOfRunOfBits(UInt32,Byte).Posit32::FractionSize().0.runningState.0\ := WaitingForStarted;
                            \Posit32::FractionSize().0.Posit32::LengthOfRunOfBits(UInt32,Byte)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    


    
    
    \Posit32::GetTwosComplement(UInt32).0._Started\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32)._Started.0\;
    \Posit32::GetTwosComplement(UInt32).0.bits.parameter.In\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32).bits.parameter.Out.0\;
    \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32)._Finished.0\ <= \Posit32::GetTwosComplement(UInt32).0._Finished\;
    \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::GetTwosComplement(UInt32).return.0\ <= \Posit32::GetTwosComplement(UInt32).0.return\;
    


    
    
    \Posit32::SetZero(UInt32,UInt16).0._Started\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::SetZero(UInt32,UInt16)._Started.0\;
    \Posit32::SetZero(UInt32,UInt16).0.bits.parameter.In\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::SetZero(UInt32,UInt16).bits.parameter.Out.0\;
    \Posit32::SetZero(UInt32,UInt16).0.index.parameter.In\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::SetZero(UInt32,UInt16).index.parameter.Out.0\;
    \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::SetZero(UInt32,UInt16)._Finished.0\ <= \Posit32::SetZero(UInt32,UInt16).0._Finished\;
    \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.Posit32::SetZero(UInt32,UInt16).return.0\ <= \Posit32::SetZero(UInt32,UInt16).0.return\;
    


    
    
    \Posit32::GetRegimeKValue().0._Started\ <= \Posit32::CalculateScaleFactor().0.Posit32::GetRegimeKValue()._Started.0\;
    \Posit32::GetRegimeKValue().0.this.parameter.In\ <= \Posit32::CalculateScaleFactor().0.Posit32::GetRegimeKValue().this.parameter.Out.0\;
    \Posit32::CalculateScaleFactor().0.Posit32::GetRegimeKValue()._Finished.0\ <= \Posit32::GetRegimeKValue().0._Finished\;
    \Posit32::CalculateScaleFactor().0.Posit32::GetRegimeKValue().return.0\ <= \Posit32::GetRegimeKValue().0.return\;
    


    
    
    \Posit32::GetExponentValue().0._Started\ <= \Posit32::CalculateScaleFactor().0.Posit32::GetExponentValue()._Started.0\;
    \Posit32::GetExponentValue().0.this.parameter.In\ <= \Posit32::CalculateScaleFactor().0.Posit32::GetExponentValue().this.parameter.Out.0\;
    \Posit32::CalculateScaleFactor().0.Posit32::GetExponentValue()._Finished.0\ <= \Posit32::GetExponentValue().0._Finished\;
    \Posit32::CalculateScaleFactor().0.Posit32::GetExponentValue().return.0\ <= \Posit32::GetExponentValue().0.return\;
    


    
    
    \Posit32::ExponentSize().0._Started\ <= \Posit32::GetExponentValue().0.Posit32::ExponentSize()._Started.0\;
    \Posit32::ExponentSize().0.this.parameter.In\ <= \Posit32::GetExponentValue().0.Posit32::ExponentSize().this.parameter.Out.0\;
    \Posit32::GetExponentValue().0.Posit32::ExponentSize()._Finished.0\ <= \Posit32::ExponentSize().0._Finished\;
    \Posit32::GetExponentValue().0.Posit32::ExponentSize().return.0\ <= \Posit32::ExponentSize().0.return\;
    


    
    \Hast::InternalInvocationProxy().Posit32::FractionSize()\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Posit32::FractionSize().Posit32::GetExponentValue().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Posit32::FractionSize().Posit32::GetExponentValue().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Posit32::FractionSize().Posit32::FractionWithHiddenBit().0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Posit32::FractionSize().Posit32::FractionWithHiddenBit().0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Posit32::FractionSize().Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Posit32::FractionSize().Quire Posit32::op_Explicit(Posit32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Hast::InternalInvocationProxy().Posit32::FractionSize().Posit32::GetExponentValue().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Posit32::FractionSize().Posit32::GetExponentValue().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Posit32::FractionSize().Posit32::FractionWithHiddenBit().0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Posit32::FractionSize().Posit32::FractionWithHiddenBit().0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Posit32::FractionSize().Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Posit32::FractionSize().Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForStarted;
                \Posit32::GetExponentValue().0.Posit32::FractionSize()._Finished.0\ <= false;
                \Posit32::FractionWithHiddenBit().0.Posit32::FractionSize()._Finished.0\ <= false;
                \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionSize()._Finished.0\ <= false;
            else 

                
                case \Hast::InternalInvocationProxy().Posit32::FractionSize().Posit32::GetExponentValue().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Posit32::GetExponentValue().0.Posit32::FractionSize()._Started.0\) then 
                            \Posit32::GetExponentValue().0.Posit32::FractionSize()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Posit32::FractionSize().Posit32::GetExponentValue().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Posit32::FractionSize().Posit32::GetExponentValue().0.runningIndex.0\ := 0;
                            \Posit32::FractionSize().0._Started\ <= true;
                            \Posit32::FractionSize().0.this.parameter.In\ <= \Posit32::GetExponentValue().0.Posit32::FractionSize().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Posit32::FractionSize().Posit32::GetExponentValue().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Posit32::FractionSize().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Posit32::FractionSize().Posit32::GetExponentValue().0.runningState.0\ := AfterFinished;
                                    \Posit32::GetExponentValue().0.Posit32::FractionSize()._Finished.0\ <= true;
                                    \Posit32::FractionSize().0._Started\ <= false;
                                    \Posit32::GetExponentValue().0.Posit32::FractionSize().return.0\ <= \Posit32::FractionSize().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Posit32::GetExponentValue().0.Posit32::FractionSize()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Posit32::FractionSize().Posit32::GetExponentValue().0.runningState.0\ := WaitingForStarted;
                            \Posit32::GetExponentValue().0.Posit32::FractionSize()._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Posit32::FractionSize().Posit32::FractionWithHiddenBit().0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Posit32::FractionWithHiddenBit().0.Posit32::FractionSize()._Started.0\) then 
                            \Posit32::FractionWithHiddenBit().0.Posit32::FractionSize()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Posit32::FractionSize().Posit32::FractionWithHiddenBit().0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Posit32::FractionSize().Posit32::FractionWithHiddenBit().0.runningIndex.0\ := 0;
                            \Posit32::FractionSize().0._Started\ <= true;
                            \Posit32::FractionSize().0.this.parameter.In\ <= \Posit32::FractionWithHiddenBit().0.Posit32::FractionSize().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Posit32::FractionSize().Posit32::FractionWithHiddenBit().0.runningIndex.0\ is 
                            when 0 => 
                                if (\Posit32::FractionSize().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Posit32::FractionSize().Posit32::FractionWithHiddenBit().0.runningState.0\ := AfterFinished;
                                    \Posit32::FractionWithHiddenBit().0.Posit32::FractionSize()._Finished.0\ <= true;
                                    \Posit32::FractionSize().0._Started\ <= false;
                                    \Posit32::FractionWithHiddenBit().0.Posit32::FractionSize().return.0\ <= \Posit32::FractionSize().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Posit32::FractionWithHiddenBit().0.Posit32::FractionSize()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Posit32::FractionSize().Posit32::FractionWithHiddenBit().0.runningState.0\ := WaitingForStarted;
                            \Posit32::FractionWithHiddenBit().0.Posit32::FractionSize()._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Posit32::FractionSize().Quire Posit32::op_Explicit(Posit32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionSize()._Started.0\) then 
                            \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionSize()._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Posit32::FractionSize().Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Posit32::FractionSize().Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ := 0;
                            \Posit32::FractionSize().0._Started\ <= true;
                            \Posit32::FractionSize().0.this.parameter.In\ <= \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionSize().this.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Posit32::FractionSize().Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Posit32::FractionSize().0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Posit32::FractionSize().Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := AfterFinished;
                                    \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionSize()._Finished.0\ <= true;
                                    \Posit32::FractionSize().0._Started\ <= false;
                                    \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionSize().return.0\ <= \Posit32::FractionSize().0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionSize()._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Posit32::FractionSize().Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForStarted;
                            \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionSize()._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    


    
    
    \Posit32::SetOne(UInt32,UInt16).0._Started\ <= \Posit32::FractionWithHiddenBit().0.Posit32::SetOne(UInt32,UInt16)._Started.0\;
    \Posit32::SetOne(UInt32,UInt16).0.this.parameter.In\ <= \Posit32::FractionWithHiddenBit().0.Posit32::SetOne(UInt32,UInt16).this.parameter.Out.0\;
    \Posit32::SetOne(UInt32,UInt16).0.bits.parameter.In\ <= \Posit32::FractionWithHiddenBit().0.Posit32::SetOne(UInt32,UInt16).bits.parameter.Out.0\;
    \Posit32::SetOne(UInt32,UInt16).0.index.parameter.In\ <= \Posit32::FractionWithHiddenBit().0.Posit32::SetOne(UInt32,UInt16).index.parameter.Out.0\;
    \Posit32::FractionWithHiddenBit().0.Posit32::SetOne(UInt32,UInt16)._Finished.0\ <= \Posit32::SetOne(UInt32,UInt16).0._Finished\;
    \Posit32::FractionWithHiddenBit().0.Posit32::SetOne(UInt32,UInt16).return.0\ <= \Posit32::SetOne(UInt32,UInt16).0.return\;
    


    
    \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Quire::op_Addition(Quire,UInt32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Quire::op_Addition(Quire,UInt32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\ := WaitingForStarted;
                \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Finished.0\ <= false;
                \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Finished.0\ <= false;
            else 

                
                case \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Started.0\) then 
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ := 0;
                            \Quire::.ctor(UInt32,UInt16).0._Started\ <= true;
                            \Quire::.ctor(UInt32,UInt16).0.this.parameter.In\ <= \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).this.parameter.Out.0\;
                            \Quire::.ctor(UInt32,UInt16).0.firstSegment.parameter.In\ <= \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).firstSegment.parameter.Out.0\;
                            \Quire::.ctor(UInt32,UInt16).0.size.parameter.In\ <= \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire::.ctor(UInt32,UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := AfterFinished;
                                    \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Finished.0\ <= true;
                                    \Quire::.ctor(UInt32,UInt16).0._Started\ <= false;
                                    \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).this.parameter.In.0\ <= \Quire::.ctor(UInt32,UInt16).0.this.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForStarted;
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Started.0\) then 
                            \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Quire::op_Addition(Quire,UInt32).0.runningIndex.0\ := 0;
                            \Quire::.ctor(UInt32,UInt16).0._Started\ <= true;
                            \Quire::.ctor(UInt32,UInt16).0.this.parameter.In\ <= \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).this.parameter.Out.0\;
                            \Quire::.ctor(UInt32,UInt16).0.firstSegment.parameter.In\ <= \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).firstSegment.parameter.Out.0\;
                            \Quire::.ctor(UInt32,UInt16).0.size.parameter.In\ <= \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Quire::op_Addition(Quire,UInt32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire::.ctor(UInt32,UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\ := AfterFinished;
                                    \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Finished.0\ <= true;
                                    \Quire::.ctor(UInt32,UInt16).0._Started\ <= false;
                                    \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).this.parameter.In.0\ <= \Quire::.ctor(UInt32,UInt16).0.this.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\ := WaitingForStarted;
                            \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    


    
    
    \Boolean Quire::op_Equality(Quire,Quire).0._Started\ <= \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire)._Started.0\;
    \Boolean Quire::op_Equality(Quire,Quire).0.left.parameter.In\ <= \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).left.parameter.Out.0\;
    \Boolean Quire::op_Equality(Quire,Quire).0.right.parameter.In\ <= \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).right.parameter.Out.0\;
    \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire)._Finished.0\ <= \Boolean Quire::op_Equality(Quire,Quire).0._Finished\;
    \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).return.0\ <= \Boolean Quire::op_Equality(Quire,Quire).0.return\;
    \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).left.parameter.In.0\ <= \Boolean Quire::op_Equality(Quire,Quire).0.left.parameter.Out\;
    \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).right.parameter.In.0\ <= \Boolean Quire::op_Equality(Quire,Quire).0.right.parameter.Out\;
    


    
    
    \Posit32::IsNaN().0._Started\ <= \Posit32::FusedSum(Posit32[],Quire).0.Posit32::IsNaN()._Started.0\;
    \Posit32::IsNaN().0.this.parameter.In\ <= \Posit32::FusedSum(Posit32[],Quire).0.Posit32::IsNaN().this.parameter.Out.0\;
    \Posit32::FusedSum(Posit32[],Quire).0.Posit32::IsNaN()._Finished.0\ <= \Posit32::IsNaN().0._Finished\;
    \Posit32::FusedSum(Posit32[],Quire).0.Posit32::IsNaN().return.0\ <= \Posit32::IsNaN().0.return\;
    


    
    \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Quire Quire::op_Addition(Quire,UInt32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Quire Quire::op_Addition(Quire,UInt32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\ := WaitingForStarted;
                \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\ <= false;
                \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\ <= false;
            else 

                
                case \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\) then 
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ := 0;
                            \Quire Quire::op_Addition(Quire,Quire).0._Started\ <= true;
                            \Quire Quire::op_Addition(Quire,Quire).0.left.parameter.In\ <= \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.Out.0\;
                            \Quire Quire::op_Addition(Quire,Quire).0.right.parameter.In\ <= \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire Quire::op_Addition(Quire,Quire).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := AfterFinished;
                                    \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\ <= true;
                                    \Quire Quire::op_Addition(Quire,Quire).0._Started\ <= false;
                                    \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).return.0\ <= \Quire Quire::op_Addition(Quire,Quire).0.return\;
                                    \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.In.0\ <= \Quire Quire::op_Addition(Quire,Quire).0.left.parameter.Out\;
                                    \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.In.0\ <= \Quire Quire::op_Addition(Quire,Quire).0.right.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForStarted;
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\) then 
                            \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Quire Quire::op_Addition(Quire,UInt32).0.runningIndex.0\ := 0;
                            \Quire Quire::op_Addition(Quire,Quire).0._Started\ <= true;
                            \Quire Quire::op_Addition(Quire,Quire).0.left.parameter.In\ <= \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.Out.0\;
                            \Quire Quire::op_Addition(Quire,Quire).0.right.parameter.In\ <= \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Quire Quire::op_Addition(Quire,UInt32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire Quire::op_Addition(Quire,Quire).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\ := AfterFinished;
                                    \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\ <= true;
                                    \Quire Quire::op_Addition(Quire,Quire).0._Started\ <= false;
                                    \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).return.0\ <= \Quire Quire::op_Addition(Quire,Quire).0.return\;
                                    \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.In.0\ <= \Quire Quire::op_Addition(Quire,Quire).0.left.parameter.Out\;
                                    \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.In.0\ <= \Quire Quire::op_Addition(Quire,Quire).0.right.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\ := WaitingForStarted;
                            \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    


    
    
    \Posit32::FractionWithHiddenBit().0._Started\ <= \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionWithHiddenBit()._Started.0\;
    \Posit32::FractionWithHiddenBit().0.this.parameter.In\ <= \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionWithHiddenBit().this.parameter.Out.0\;
    \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionWithHiddenBit()._Finished.0\ <= \Posit32::FractionWithHiddenBit().0._Finished\;
    \Quire Posit32::op_Explicit(Posit32).0.Posit32::FractionWithHiddenBit().return.0\ <= \Posit32::FractionWithHiddenBit().0.return\;
    


    
    \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Posit32::op_Explicit(Posit32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_Addition(Quire,Quire).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_Addition(Quire,Quire).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_RightShift(Quire,Int32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_RightShift(Quire,Int32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_LeftShift(Quire,Int32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_LeftShift(Quire,Int32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_Addition(Quire,Quire).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_Addition(Quire,Quire).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_RightShift(Quire,Int32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_RightShift(Quire,Int32).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_LeftShift(Quire,Int32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_LeftShift(Quire,Int32).0.runningState.0\ := WaitingForStarted;
                \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
                \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
                \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
                \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
            else 

                
                case \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\) then 
                            \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ := 0;
                            \Quire::.ctor(UInt64[],UInt16).0._Started\ <= true;
                            \Quire::.ctor(UInt64[],UInt16).0.this.parameter.In\ <= \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\;
                            \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.In\ <= \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\;
                            \Quire::.ctor(UInt64[],UInt16).0.size.parameter.In\ <= \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire::.ctor(UInt64[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := AfterFinished;
                                    \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= true;
                                    \Quire::.ctor(UInt64[],UInt16).0._Started\ <= false;
                                    \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\ <= \Quire::.ctor(UInt64[],UInt16).0.this.parameter.Out\;
                                    \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\ <= \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForStarted;
                            \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_Addition(Quire,Quire).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Started.0\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_Addition(Quire,Quire).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_Addition(Quire,Quire).0.runningIndex.0\ := 0;
                            \Quire::.ctor(UInt64[],UInt16).0._Started\ <= true;
                            \Quire::.ctor(UInt64[],UInt16).0.this.parameter.In\ <= \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\;
                            \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.In\ <= \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\;
                            \Quire::.ctor(UInt64[],UInt16).0.size.parameter.In\ <= \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_Addition(Quire,Quire).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire::.ctor(UInt64[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_Addition(Quire,Quire).0.runningState.0\ := AfterFinished;
                                    \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= true;
                                    \Quire::.ctor(UInt64[],UInt16).0._Started\ <= false;
                                    \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\ <= \Quire::.ctor(UInt64[],UInt16).0.this.parameter.Out\;
                                    \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\ <= \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_Addition(Quire,Quire).0.runningState.0\ := WaitingForStarted;
                            \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_RightShift(Quire,Int32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\) then 
                            \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_RightShift(Quire,Int32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_RightShift(Quire,Int32).0.runningIndex.0\ := 0;
                            \Quire::.ctor(UInt64[],UInt16).0._Started\ <= true;
                            \Quire::.ctor(UInt64[],UInt16).0.this.parameter.In\ <= \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\;
                            \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.In\ <= \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\;
                            \Quire::.ctor(UInt64[],UInt16).0.size.parameter.In\ <= \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_RightShift(Quire,Int32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire::.ctor(UInt64[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_RightShift(Quire,Int32).0.runningState.0\ := AfterFinished;
                                    \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= true;
                                    \Quire::.ctor(UInt64[],UInt16).0._Started\ <= false;
                                    \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\ <= \Quire::.ctor(UInt64[],UInt16).0.this.parameter.Out\;
                                    \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\ <= \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_RightShift(Quire,Int32).0.runningState.0\ := WaitingForStarted;
                            \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_LeftShift(Quire,Int32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\) then 
                            \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_LeftShift(Quire,Int32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_LeftShift(Quire,Int32).0.runningIndex.0\ := 0;
                            \Quire::.ctor(UInt64[],UInt16).0._Started\ <= true;
                            \Quire::.ctor(UInt64[],UInt16).0.this.parameter.In\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\;
                            \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.In\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\;
                            \Quire::.ctor(UInt64[],UInt16).0.size.parameter.In\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_LeftShift(Quire,Int32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire::.ctor(UInt64[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_LeftShift(Quire,Int32).0.runningState.0\ := AfterFinished;
                                    \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= true;
                                    \Quire::.ctor(UInt64[],UInt16).0._Started\ <= false;
                                    \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\ <= \Quire::.ctor(UInt64[],UInt16).0.this.parameter.Out\;
                                    \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\ <= \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_LeftShift(Quire,Int32).0.runningState.0\ := WaitingForStarted;
                            \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    


    
    
    \Posit32::CalculateScaleFactor().0._Started\ <= \Quire Posit32::op_Explicit(Posit32).0.Posit32::CalculateScaleFactor()._Started.0\;
    \Posit32::CalculateScaleFactor().0.this.parameter.In\ <= \Quire Posit32::op_Explicit(Posit32).0.Posit32::CalculateScaleFactor().this.parameter.Out.0\;
    \Quire Posit32::op_Explicit(Posit32).0.Posit32::CalculateScaleFactor()._Finished.0\ <= \Posit32::CalculateScaleFactor().0._Finished\;
    \Quire Posit32::op_Explicit(Posit32).0.Posit32::CalculateScaleFactor().return.0\ <= \Posit32::CalculateScaleFactor().0.return\;
    


    
    
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._Started\ <= \Hast::ExternalInvocationProxy().Posit32FusedCalculator::CalculateFusedSum(SimpleMemory)._Started.0\;
    \Hast::ExternalInvocationProxy().Posit32FusedCalculator::CalculateFusedSum(SimpleMemory)._Finished.0\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._Finished\;
    


    
    \CellIndex\ <= to_integer(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.CellIndex\) when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.ReadEnable\ or \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.WriteEnable\ else 0;
    \DataOut\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.DataOut\ when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.WriteEnable\ else (others => '0');
    \ReadEnable\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.ReadEnable\;
    \WriteEnable\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.WriteEnable\;
    

end Imp;





library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package TypeConversion is
    function SmartResize(input: unsigned; size: natural) return unsigned;
    function SmartResize(input: signed; size: natural) return signed;
    function ToUnsignedAndExpand(input: signed; size: natural) return unsigned;
end TypeConversion;
        
package body TypeConversion is

    
    
    
    
    
    
    function SmartResize(input: unsigned; size: natural) return unsigned is
    begin
        if (size < input'LENGTH) then
            return input(size - 1 downto 0);
        else
            
            
            
            return resize(input, size);
        end if;
    end SmartResize;

    function SmartResize(input: signed; size: natural) return signed is
    begin
        if (size < input'LENGTH) then
            return input(size - 1 downto 0);
        else
            return resize(input, size);
        end if;
    end SmartResize;

    function ToUnsignedAndExpand(input: signed; size: natural) return unsigned is
        variable result: unsigned(size - 1 downto 0);
    begin
        if (input >= 0) then
            return resize(unsigned(input), size);
        else 
            result := (others => '1');
            result(input'LENGTH - 1 downto 0) := unsigned(input);
            return result;
        end if;
    end ToUnsignedAndExpand;

end TypeConversion;


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
        
package SimpleMemory is
    
    function ConvertUInt32ToStdLogicVector(input: unsigned(31 downto 0)) return std_logic_vector;
    function ConvertStdLogicVectorToUInt32(input : std_logic_vector) return unsigned;
        
    function ConvertBooleanToStdLogicVector(input: boolean) return std_logic_vector;
    function ConvertStdLogicVectorToBoolean(input : std_logic_vector) return boolean;
        
    function ConvertInt32ToStdLogicVector(input: signed(31 downto 0)) return std_logic_vector;
    function ConvertStdLogicVectorToInt32(input : std_logic_vector) return signed;
end SimpleMemory;
        
package body SimpleMemory is

    function ConvertUInt32ToStdLogicVector(input: unsigned(31 downto 0)) return std_logic_vector is
    begin
        return std_logic_vector(input);
    end ConvertUInt32ToStdLogicVector;
    
    function ConvertStdLogicVectorToUInt32(input : std_logic_vector) return unsigned is
    begin
        return unsigned(input);
    end ConvertStdLogicVectorToUInt32;
    
    function ConvertBooleanToStdLogicVector(input: boolean) return std_logic_vector is 
    begin
        case input is
            when true => return X"FFFFFFFF";
            when false => return X"00000000";
            when others => return X"00000000";
        end case;
    end ConvertBooleanToStdLogicVector;

    function ConvertStdLogicVectorToBoolean(input : std_logic_vector) return boolean is 
    begin
        
        return not(input = X"00000000");
    end ConvertStdLogicVectorToBoolean;

    function ConvertInt32ToStdLogicVector(input: signed(31 downto 0)) return std_logic_vector is
    begin
        return std_logic_vector(input);
    end ConvertInt32ToStdLogicVector;

    function ConvertStdLogicVectorToInt32(input : std_logic_vector) return signed is
    begin
        return signed(input);
    end ConvertStdLogicVectorToInt32;

end SimpleMemory;


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.TypeConversion.all;
library work;
use work.SimpleMemory.all;

entity Hast_IP is 
    port(
        \DataIn\: In std_logic_vector(31 downto 0);
        \DataOut\: Out std_logic_vector(31 downto 0);
        \CellIndex\: Out integer;
        \ReadEnable\: Out boolean;
        \WriteEnable\: Out boolean;
        \ReadsDone\: In boolean;
        \WritesDone\: In boolean;
        \MemberId\: In integer;
        \Reset\: In std_logic;
        \Started\: In boolean;
        \Finished\: Out boolean;
        \Clock\: In std_logic
    );
    
    
    

    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    

end Hast_IP;

architecture Imp of Hast_IP is 
    
    
    
    
    
    
    
    
    

    
    attribute altera_attribute: string;
    attribute altera_attribute of Imp: architecture is "-name SDC_STATEMENT ""set_multicycle_path 8 -setup -to {*Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._StateMachine:Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.0[*]}"";-name SDC_STATEMENT ""set_multicycle_path 7 -hold -to {*Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._StateMachine:Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.0[*]}"";-name SDC_STATEMENT ""set_multicycle_path 8 -setup -to {*Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._StateMachine:Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.1[*]}"";-name SDC_STATEMENT ""set_multicycle_path 7 -hold -to {*Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._StateMachine:Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.1[*]}""";


    
    type \Lombiq.Arithmetics.Posit32\ is record 
        \IsNull\: boolean;
        \PositBits\: unsigned(31 downto 0);
    end record;
    type \Lombiq.Arithmetics.Posit32_Array\ is array (integer range <>) of \Lombiq.Arithmetics.Posit32\;
    type \unsigned64_Array\ is array (integer range <>) of unsigned(63 downto 0);
    type \Lombiq.Arithmetics.Quire\ is record 
        \IsNull\: boolean;
        \Size\: unsigned(15 downto 0);
        \SegmentCount\: unsigned(15 downto 0);
        \Segments\: \unsigned64_Array\(0 to 7);
    end record;
    


    
    
    type \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._States\ is (
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_0\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_1\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_2\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_3\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_4\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_5\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_6\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_7\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_8\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_9\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_10\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_11\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_12\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_13\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_14\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_15\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_16\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_17\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_18\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_19\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_20\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_21\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_22\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_23\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_24\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_25\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_26\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_27\, 
        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_28\);
    
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._Finished\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.CellIndex\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.DataOut\: std_logic_vector(31 downto 0) := (others => '0');
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.ReadEnable\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.WriteEnable\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).this.parameter.Out.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).value.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Started.0\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32).x.parameter.Out.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Started.0\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).this.parameter.Out.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).bits.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).fromBitMask.parameter.Out.0\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean)._Started.0\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).posits.parameter.Out.0\: \Lombiq.Arithmetics.Posit32_Array\(0 to 159);
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).startingValue.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire)._Started.0\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).this.parameter.Out.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).q.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire)._Started.0\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._Started\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).this.parameter.In.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Finished.0\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32).return.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).this.parameter.In.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean)._Finished.0\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).posits.parameter.In.0\: \Lombiq.Arithmetics.Posit32_Array\(0 to 159);
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).startingValue.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire)._Finished.0\: boolean := false;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).return.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).this.parameter.In.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).q.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire)._Finished.0\: boolean := false;
    


    
    
    type \Posit32::.ctor(UInt32,Boolean).0._States\ is (
        \Posit32::.ctor(UInt32,Boolean).0._State_0\, 
        \Posit32::.ctor(UInt32,Boolean).0._State_1\, 
        \Posit32::.ctor(UInt32,Boolean).0._State_2\);
    
    Signal \Posit32::.ctor(UInt32,Boolean).0._Finished\: boolean := false;
    Signal \Posit32::.ctor(UInt32,Boolean).0.this.parameter.Out\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::.ctor(UInt32,Boolean).0._Started\: boolean := false;
    Signal \Posit32::.ctor(UInt32,Boolean).0.this.parameter.In\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::.ctor(UInt32,Boolean).0.bits.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::.ctor(UInt32,Boolean).0.fromBitMask.parameter.In\: boolean := false;
    


    
    
    type \Posit32::.ctor(Quire).0._States\ is (
        \Posit32::.ctor(Quire).0._State_0\, 
        \Posit32::.ctor(Quire).0._State_1\, 
        \Posit32::.ctor(Quire).0._State_2\, 
        \Posit32::.ctor(Quire).0._State_3\, 
        \Posit32::.ctor(Quire).0._State_4\, 
        \Posit32::.ctor(Quire).0._State_5\, 
        \Posit32::.ctor(Quire).0._State_6\, 
        \Posit32::.ctor(Quire).0._State_7\, 
        \Posit32::.ctor(Quire).0._State_8\, 
        \Posit32::.ctor(Quire).0._State_9\, 
        \Posit32::.ctor(Quire).0._State_10\, 
        \Posit32::.ctor(Quire).0._State_11\, 
        \Posit32::.ctor(Quire).0._State_12\, 
        \Posit32::.ctor(Quire).0._State_13\, 
        \Posit32::.ctor(Quire).0._State_14\, 
        \Posit32::.ctor(Quire).0._State_15\, 
        \Posit32::.ctor(Quire).0._State_16\, 
        \Posit32::.ctor(Quire).0._State_17\, 
        \Posit32::.ctor(Quire).0._State_18\, 
        \Posit32::.ctor(Quire).0._State_19\, 
        \Posit32::.ctor(Quire).0._State_20\, 
        \Posit32::.ctor(Quire).0._State_21\, 
        \Posit32::.ctor(Quire).0._State_22\, 
        \Posit32::.ctor(Quire).0._State_23\, 
        \Posit32::.ctor(Quire).0._State_24\);
    
    Signal \Posit32::.ctor(Quire).0._Finished\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.this.parameter.Out\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::.ctor(Quire).0.q.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).right.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).x.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire).q.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire)._Started.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).left.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).right.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32)._Started.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire).x.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire)._Started.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).signBit.parameter.Out.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).regimeKValue.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).exponentBits.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).fractionBits.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32)._Started.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0._Started\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.this.parameter.In\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::.ctor(Quire).0.q.parameter.In\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Finished.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).return.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).x.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Finished.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).return.0\: unsigned(63 downto 0) := to_unsigned(0, 64);
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire).q.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire)._Finished.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire).return.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).left.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32)._Finished.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).return.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).return.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire).x.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire)._Finished.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32)._Finished.0\: boolean := false;
    Signal \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).return.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    


    
    
    type \Posit32::.ctor(UInt32).0._States\ is (
        \Posit32::.ctor(UInt32).0._State_0\, 
        \Posit32::.ctor(UInt32).0._State_1\, 
        \Posit32::.ctor(UInt32).0._State_2\);
    
    Signal \Posit32::.ctor(UInt32).0._Finished\: boolean := false;
    Signal \Posit32::.ctor(UInt32).0.this.parameter.Out\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::.ctor(UInt32).0._Started\: boolean := false;
    Signal \Posit32::.ctor(UInt32).0.this.parameter.In\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::.ctor(UInt32).0.value.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    


    
    
    type \Posit32::.ctor(Int32).0._States\ is (
        \Posit32::.ctor(Int32).0._State_0\, 
        \Posit32::.ctor(Int32).0._State_1\, 
        \Posit32::.ctor(Int32).0._State_2\, 
        \Posit32::.ctor(Int32).0._State_3\);
    
    Signal \Posit32::.ctor(Int32).0._Finished\: boolean := false;
    Signal \Posit32::.ctor(Int32).0.this.parameter.Out\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32).this.parameter.Out.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32).value.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32)._Started.0\: boolean := false;
    Signal \Posit32::.ctor(Int32).0._Started\: boolean := false;
    Signal \Posit32::.ctor(Int32).0.this.parameter.In\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::.ctor(Int32).0.value.parameter.In\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32).this.parameter.In.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32)._Finished.0\: boolean := false;
    


    
    
    type \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._States\ is (
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_0\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_1\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_2\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_3\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_4\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_5\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_6\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_7\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_8\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_9\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_10\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_11\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_12\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_13\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_14\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_15\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_16\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_17\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_18\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_19\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_20\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_21\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_22\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_23\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_24\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_25\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_26\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_27\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_28\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_29\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_30\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_31\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_32\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_33\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_34\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_35\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_36\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_37\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_38\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_39\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_40\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_41\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_42\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_43\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_44\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_45\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_46\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_47\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_48\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_49\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_50\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_51\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_52\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_53\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_54\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_55\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_56\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_57\, 
        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_58\);
    
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._Finished\: boolean := false;
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._Started\: boolean := false;
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.signBit.parameter.In\: boolean := false;
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.regimeKValue.parameter.In\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    


    
    
    type \Posit32::FusedSum(Posit32[],Quire).0._States\ is (
        \Posit32::FusedSum(Posit32[],Quire).0._State_0\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_1\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_2\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_3\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_4\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_5\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_6\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_7\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_8\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_9\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_10\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_11\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_12\, 
        \Posit32::FusedSum(Posit32[],Quire).0._State_13\);
    
    Signal \Posit32::FusedSum(Posit32[],Quire).0._Finished\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.return\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.posits.parameter.Out\: \Lombiq.Arithmetics.Posit32_Array\(0 to 159);
    Signal \Posit32::FusedSum(Posit32[],Quire).0.startingValue.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).this.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).firstSegment.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Started.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).left.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).right.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire)._Started.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32).x.parameter.Out.0\: \Lombiq.Arithmetics.Posit32\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Started.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0._Started\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.posits.parameter.In\: \Lombiq.Arithmetics.Posit32_Array\(0 to 159);
    Signal \Posit32::FusedSum(Posit32[],Quire).0.startingValue.parameter.In\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).this.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Finished.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).return.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).left.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).right.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire)._Finished.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).return.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32).return.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\: boolean := false;
    Signal \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).return.0\: \Lombiq.Arithmetics.Quire\;
    


    
    
    type \Quire Posit32::op_Explicit(Posit32).0._States\ is (
        \Quire Posit32::op_Explicit(Posit32).0._State_0\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_1\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_2\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_3\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_4\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_5\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_6\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_7\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_8\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_9\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_10\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_11\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_12\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_13\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_14\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_15\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_16\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_17\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_18\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_19\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_20\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_21\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_22\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_23\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_24\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_25\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_26\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_27\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_28\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_29\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_30\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_31\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_32\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_33\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_34\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_35\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_36\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_37\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_38\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_39\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_40\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_41\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_42\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_43\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_44\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_45\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_46\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_47\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_48\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_49\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_50\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_51\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_52\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_53\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_54\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_55\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_56\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_57\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_58\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_59\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_60\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_61\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_62\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_63\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_64\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_65\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_66\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_67\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_68\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_69\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_70\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_71\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_72\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_73\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_74\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_75\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_76\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_77\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_78\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_79\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_80\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_81\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_82\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_83\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_84\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_85\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_86\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_87\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_88\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_89\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_90\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_91\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_92\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_93\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_94\, 
        \Quire Posit32::op_Explicit(Posit32).0._State_95\);
    
    Signal \Quire Posit32::op_Explicit(Posit32).0._Finished\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0.return\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16).this.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16).firstSegment.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16)._Started.0\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_OnesComplement(Quire).q.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_OnesComplement(Quire)._Started.0\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32).left.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32).right.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32)._Started.0\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0._Started\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0.x.parameter.In\: \Lombiq.Arithmetics.Posit32\;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16).this.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16)._Finished.0\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).return.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_OnesComplement(Quire).q.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_OnesComplement(Quire)._Finished.0\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_OnesComplement(Quire).return.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32).left.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32)._Finished.0\: boolean := false;
    Signal \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32).return.0\: \Lombiq.Arithmetics.Quire\;
    


    
    
    type \Quire::.ctor(UInt64[],UInt16).0._States\ is (
        \Quire::.ctor(UInt64[],UInt16).0._State_0\, 
        \Quire::.ctor(UInt64[],UInt16).0._State_1\, 
        \Quire::.ctor(UInt64[],UInt16).0._State_2\, 
        \Quire::.ctor(UInt64[],UInt16).0._State_3\, 
        \Quire::.ctor(UInt64[],UInt16).0._State_4\);
    
    Signal \Quire::.ctor(UInt64[],UInt16).0._Finished\: boolean := false;
    Signal \Quire::.ctor(UInt64[],UInt16).0.this.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.Out\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
    Signal \Quire::.ctor(UInt64[],UInt16).0._Started\: boolean := false;
    Signal \Quire::.ctor(UInt64[],UInt16).0.this.parameter.In\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.In\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
    Signal \Quire::.ctor(UInt64[],UInt16).0.size.parameter.In\: unsigned(15 downto 0) := to_unsigned(0, 16);
    


    
    
    type \Quire::.ctor(UInt32,UInt16).0._States\ is (
        \Quire::.ctor(UInt32,UInt16).0._State_0\, 
        \Quire::.ctor(UInt32,UInt16).0._State_1\, 
        \Quire::.ctor(UInt32,UInt16).0._State_2\, 
        \Quire::.ctor(UInt32,UInt16).0._State_3\, 
        \Quire::.ctor(UInt32,UInt16).0._State_4\, 
        \Quire::.ctor(UInt32,UInt16).0._State_5\, 
        \Quire::.ctor(UInt32,UInt16).0._State_6\, 
        \Quire::.ctor(UInt32,UInt16).0._State_7\, 
        \Quire::.ctor(UInt32,UInt16).0._State_8\);
    
    Signal \Quire::.ctor(UInt32,UInt16).0._Finished\: boolean := false;
    Signal \Quire::.ctor(UInt32,UInt16).0.this.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire::.ctor(UInt32,UInt16).0._Started\: boolean := false;
    Signal \Quire::.ctor(UInt32,UInt16).0.this.parameter.In\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire::.ctor(UInt32,UInt16).0.firstSegment.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Quire::.ctor(UInt32,UInt16).0.size.parameter.In\: unsigned(15 downto 0) := to_unsigned(0, 16);
    


    
    
    type \Quire Quire::op_Addition(Quire,Quire).0._States\ is (
        \Quire Quire::op_Addition(Quire,Quire).0._State_0\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_1\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_2\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_3\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_4\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_5\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_6\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_7\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_8\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_9\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_10\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_11\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_12\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_13\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_14\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_15\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_16\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_17\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_18\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_19\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_20\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_21\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_22\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_23\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_24\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_25\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_26\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_27\, 
        \Quire Quire::op_Addition(Quire,Quire).0._State_28\);
    
    Signal \Quire Quire::op_Addition(Quire,Quire).0._Finished\: boolean := false;
    Signal \Quire Quire::op_Addition(Quire,Quire).0.return\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,Quire).0.left.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,Quire).0.right.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
    Signal \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Started.0\: boolean := false;
    Signal \Quire Quire::op_Addition(Quire,Quire).0._Started\: boolean := false;
    Signal \Quire Quire::op_Addition(Quire,Quire).0.left.parameter.In\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,Quire).0.right.parameter.In\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
    Signal \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\: boolean := false;
    


    
    
    type \Quire Quire::op_Addition(Quire,UInt32).0._States\ is (
        \Quire Quire::op_Addition(Quire,UInt32).0._State_0\, 
        \Quire Quire::op_Addition(Quire,UInt32).0._State_1\, 
        \Quire Quire::op_Addition(Quire,UInt32).0._State_2\, 
        \Quire Quire::op_Addition(Quire,UInt32).0._State_3\, 
        \Quire Quire::op_Addition(Quire,UInt32).0._State_4\);
    
    Signal \Quire Quire::op_Addition(Quire,UInt32).0._Finished\: boolean := false;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.return\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.left.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).this.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).firstSegment.parameter.Out.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Started.0\: boolean := false;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\: boolean := false;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0._Started\: boolean := false;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.left.parameter.In\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.right.parameter.In\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).this.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Finished.0\: boolean := false;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\: boolean := false;
    Signal \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).return.0\: \Lombiq.Arithmetics.Quire\;
    


    
    
    type \Quire Quire::op_OnesComplement(Quire).0._States\ is (
        \Quire Quire::op_OnesComplement(Quire).0._State_0\, 
        \Quire Quire::op_OnesComplement(Quire).0._State_1\, 
        \Quire Quire::op_OnesComplement(Quire).0._State_2\, 
        \Quire Quire::op_OnesComplement(Quire).0._State_3\, 
        \Quire Quire::op_OnesComplement(Quire).0._State_4\, 
        \Quire Quire::op_OnesComplement(Quire).0._State_5\);
    
    Signal \Quire Quire::op_OnesComplement(Quire).0._Finished\: boolean := false;
    Signal \Quire Quire::op_OnesComplement(Quire).0.return\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_OnesComplement(Quire).0.q.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_OnesComplement(Quire).0._Started\: boolean := false;
    Signal \Quire Quire::op_OnesComplement(Quire).0.q.parameter.In\: \Lombiq.Arithmetics.Quire\;
    


    
    
    type \Boolean Quire::op_Equality(Quire,Quire).0._States\ is (
        \Boolean Quire::op_Equality(Quire,Quire).0._State_0\, 
        \Boolean Quire::op_Equality(Quire,Quire).0._State_1\, 
        \Boolean Quire::op_Equality(Quire,Quire).0._State_2\, 
        \Boolean Quire::op_Equality(Quire,Quire).0._State_3\, 
        \Boolean Quire::op_Equality(Quire,Quire).0._State_4\, 
        \Boolean Quire::op_Equality(Quire,Quire).0._State_5\, 
        \Boolean Quire::op_Equality(Quire,Quire).0._State_6\, 
        \Boolean Quire::op_Equality(Quire,Quire).0._State_7\, 
        \Boolean Quire::op_Equality(Quire,Quire).0._State_8\);
    
    Signal \Boolean Quire::op_Equality(Quire,Quire).0._Finished\: boolean := false;
    Signal \Boolean Quire::op_Equality(Quire,Quire).0.return\: boolean := false;
    Signal \Boolean Quire::op_Equality(Quire,Quire).0.left.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Boolean Quire::op_Equality(Quire,Quire).0.right.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Boolean Quire::op_Equality(Quire,Quire).0._Started\: boolean := false;
    Signal \Boolean Quire::op_Equality(Quire,Quire).0.left.parameter.In\: \Lombiq.Arithmetics.Quire\;
    Signal \Boolean Quire::op_Equality(Quire,Quire).0.right.parameter.In\: \Lombiq.Arithmetics.Quire\;
    


    
    
    type \Quire Quire::op_RightShift(Quire,Int32).0._States\ is (
        \Quire Quire::op_RightShift(Quire,Int32).0._State_0\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_1\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_2\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_3\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_4\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_5\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_6\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_7\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_8\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_9\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_10\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_11\, 
        \Quire Quire::op_RightShift(Quire,Int32).0._State_12\);
    
    Signal \Quire Quire::op_RightShift(Quire,Int32).0._Finished\: boolean := false;
    Signal \Quire Quire::op_RightShift(Quire,Int32).0.return\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_RightShift(Quire,Int32).0.left.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
    Signal \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\: boolean := false;
    Signal \Quire Quire::op_RightShift(Quire,Int32).0._Started\: boolean := false;
    Signal \Quire Quire::op_RightShift(Quire,Int32).0.left.parameter.In\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_RightShift(Quire,Int32).0.right.parameter.In\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
    Signal \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\: boolean := false;
    


    
    
    type \Quire Quire::op_LeftShift(Quire,Int32).0._States\ is (
        \Quire Quire::op_LeftShift(Quire,Int32).0._State_0\, 
        \Quire Quire::op_LeftShift(Quire,Int32).0._State_1\, 
        \Quire Quire::op_LeftShift(Quire,Int32).0._State_2\, 
        \Quire Quire::op_LeftShift(Quire,Int32).0._State_3\, 
        \Quire Quire::op_LeftShift(Quire,Int32).0._State_4\, 
        \Quire Quire::op_LeftShift(Quire,Int32).0._State_5\, 
        \Quire Quire::op_LeftShift(Quire,Int32).0._State_6\, 
        \Quire Quire::op_LeftShift(Quire,Int32).0._State_7\, 
        \Quire Quire::op_LeftShift(Quire,Int32).0._State_8\, 
        \Quire Quire::op_LeftShift(Quire,Int32).0._State_9\, 
        \Quire Quire::op_LeftShift(Quire,Int32).0._State_10\);
    
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0._Finished\: boolean := false;
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0.return\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0.left.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\: boolean := false;
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0._Started\: boolean := false;
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0.left.parameter.In\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0.right.parameter.In\: signed(31 downto 0) := to_signed(0, 32);
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\: \Lombiq.Arithmetics.Quire\;
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
    Signal \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\: boolean := false;
    


    
    
    type \UInt64 Quire::op_Explicit(Quire).0._States\ is (
        \UInt64 Quire::op_Explicit(Quire).0._State_0\, 
        \UInt64 Quire::op_Explicit(Quire).0._State_1\, 
        \UInt64 Quire::op_Explicit(Quire).0._State_2\);
    
    Signal \UInt64 Quire::op_Explicit(Quire).0._Finished\: boolean := false;
    Signal \UInt64 Quire::op_Explicit(Quire).0.return\: unsigned(63 downto 0) := to_unsigned(0, 64);
    Signal \UInt64 Quire::op_Explicit(Quire).0.x.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \UInt64 Quire::op_Explicit(Quire).0._Started\: boolean := false;
    Signal \UInt64 Quire::op_Explicit(Quire).0.x.parameter.In\: \Lombiq.Arithmetics.Quire\;
    


    
    
    type \UInt32 Quire::op_Explicit(Quire).0._States\ is (
        \UInt32 Quire::op_Explicit(Quire).0._State_0\, 
        \UInt32 Quire::op_Explicit(Quire).0._State_1\, 
        \UInt32 Quire::op_Explicit(Quire).0._State_2\);
    
    Signal \UInt32 Quire::op_Explicit(Quire).0._Finished\: boolean := false;
    Signal \UInt32 Quire::op_Explicit(Quire).0.return\: unsigned(31 downto 0) := to_unsigned(0, 32);
    Signal \UInt32 Quire::op_Explicit(Quire).0.x.parameter.Out\: \Lombiq.Arithmetics.Quire\;
    Signal \UInt32 Quire::op_Explicit(Quire).0._Started\: boolean := false;
    Signal \UInt32 Quire::op_Explicit(Quire).0.x.parameter.In\: \Lombiq.Arithmetics.Quire\;
    


    
    
    Signal \FinishedInternal\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().Posit32FusedCalculator::CalculateFusedSum(SimpleMemory)._Started.0\: boolean := false;
    Signal \Hast::ExternalInvocationProxy().Posit32FusedCalculator::CalculateFusedSum(SimpleMemory)._Finished.0\: boolean := false;
    


    
    type \InternalInvocationProxy_boolean_Array\ is array (integer range <>) of boolean;
    type \Hast::InternalInvocationProxy()._RunningStates\ is (
        WaitingForStarted, 
        WaitingForFinished, 
        AfterFinished);
    

begin 

    
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._StateMachine\: process (\Clock\) 
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\: \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._States\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_0\;
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.dataIn.0\: std_logic_vector(31 downto 0) := (others => '0');
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.array\: \Lombiq.Arithmetics.Posit32_Array\(0 to 159);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.quire\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectde41e31d213f26bcb14dc4059ca0ea22b32147dbfb27f3d69d5ff482204eea98\: \Lombiq.Arithmetics.Posit32\;
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.return.0\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.3\: signed(63 downto 0) := to_signed(0, 64);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.4\: boolean := false;
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.5\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num3\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.6\: boolean := false;
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.7\: boolean := false;
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.8\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.9\: signed(63 downto 0) := to_signed(0, 64);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.10\: boolean := false;
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.11\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.12\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.13\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.dataIn.1\: std_logic_vector(31 downto 0) := (others => '0');
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.14\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.return.1\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.15\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectffd9139c321969eb0a42e1e3ae043fc0d22d96a54e32c2dc05d540c7e97af68e\: \Lombiq.Arithmetics.Posit32\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._Finished\ <= false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.DataOut\ <= (others => '0');
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).value.parameter.Out.0\ <= to_signed(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Started.0\ <= false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Started.0\ <= false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).bits.parameter.Out.0\ <= to_unsigned(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).fromBitMask.parameter.Out.0\ <= false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean)._Started.0\ <= false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire)._Started.0\ <= false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire)._Started.0\ <= false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_0\;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num\ := to_unsigned(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.dataIn.0\ := (others => '0');
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num2\ := to_unsigned(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.0\ := to_unsigned(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.1\ := to_unsigned(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.1\ := to_signed(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.2\ := to_unsigned(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.3\ := to_signed(0, 64);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.4\ := false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.5\ := to_unsigned(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num3\ := to_signed(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.6\ := false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\ := to_signed(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.7\ := false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.8\ := to_signed(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.9\ := to_signed(0, 64);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.10\ := false;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.11\ := to_signed(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.12\ := to_signed(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.13\ := to_signed(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.dataIn.1\ := (others => '0');
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.14\ := to_signed(0, 32);
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.15\ := to_signed(0, 32);
            else 
                case \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ is 
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_0\ => 
                        
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._Started\ = true) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_2\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_1\ => 
                        
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._Started\ = true) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._Finished\ <= true;
                        else 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._Finished\ <= false;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_0\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_2\ => 
                        
                        
                        
                        
                        
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.ReadEnable\ <= true;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_3\;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_3\ => 
                        
                        if (\ReadsDone\ = true) then 
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.dataIn.0\ := \DataIn\;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num\ := ConvertStdLogicVectorToUInt32(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.dataIn.0\);
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectde41e31d213f26bcb14dc4059ca0ea22b32147dbfb27f3d69d5ff482204eea98\.\IsNull\ := false;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectde41e31d213f26bcb14dc4059ca0ea22b32147dbfb27f3d69d5ff482204eea98\.\PositBits\ := to_unsigned(0, 32);
                            
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).this.parameter.Out.0\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectde41e31d213f26bcb14dc4059ca0ea22b32147dbfb27f3d69d5ff482204eea98\;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).value.parameter.Out.0\ <= to_signed(0, 32);
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Started.0\ <= true;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_4\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_4\ => 
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Started.0\ = \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Finished.0\) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Started.0\ <= false;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectde41e31d213f26bcb14dc4059ca0ea22b32147dbfb27f3d69d5ff482204eea98\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).this.parameter.In.0\;
                            
                            
                            
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32).x.parameter.Out.0\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectde41e31d213f26bcb14dc4059ca0ea22b32147dbfb27f3d69d5ff482204eea98\;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Started.0\ <= true;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_5\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_5\ => 
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Started.0\ = \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Started.0\ <= false;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.return.0\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32).return.0\;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.quire\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.return.0\;
                            
                            
                            
                            
                            
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_6\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_6\ => 
                        
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.0\ >= to_signed(8, 32)) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_7\;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.0\ := to_signed(0, 32);
                        else 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.0\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.0\ + to_signed(1, 32);
                        end if;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.0\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num\ / to_unsigned(160, 32);
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_7\ => 
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num2\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.0\;
                        
                        
                        
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_8\;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_8\ => 
                        
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.1\ >= to_signed(8, 32)) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_9\;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.1\ := to_signed(0, 32);
                        else 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.1\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.clockCyclesWaitedForBinaryOperationResult.1\ + to_signed(1, 32);
                        end if;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.1\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num\ / to_unsigned(160, 32);
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_9\ => 
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.2\ := SmartResize(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.1\ * to_unsigned(160, 32), 32);
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.3\ := signed(SmartResize(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num\ - \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.2\, 64));
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_10\;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_10\ => 
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.4\ := (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.3\) /= to_signed(0, 64);

                        
                        
                        

                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.4\) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_12\;
                        else 
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_11\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_11\ => 
                        
                        
                        
                        
                        
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num3\ := to_signed(0, 32);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_13\;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_12\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.5\ := SmartResize(unsigned(signed(SmartResize((\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num2\), 64)) + to_signed(1, 64)), 32);
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num2\ := (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.5\);
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ = \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_12\) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_11\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_13\ => 
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.6\ := SmartResize((\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num3\), 64) < signed(SmartResize((\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num2\), 64));
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.6\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\ := to_signed(0, 32);
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_15\;
                        else 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_14\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_14\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectffd9139c321969eb0a42e1e3ae043fc0d22d96a54e32c2dc05d540c7e97af68e\.\IsNull\ := false;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectffd9139c321969eb0a42e1e3ae043fc0d22d96a54e32c2dc05d540c7e97af68e\.\PositBits\ := to_unsigned(0, 32);
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).this.parameter.Out.0\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectffd9139c321969eb0a42e1e3ae043fc0d22d96a54e32c2dc05d540c7e97af68e\;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).q.parameter.Out.0\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.quire\;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire)._Started.0\ <= true;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_27\;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_15\ => 
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.7\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\ < to_signed(160, 32);
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.7\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.8\ := SmartResize(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num3\ * to_signed(160, 32), 32);
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_17\;
                        else 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_16\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_16\ => 
                        
                        
                        
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).posits.parameter.Out.0\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.array\;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).startingValue.parameter.Out.0\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.quire\;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire)._Started.0\ <= true;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_26\;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_17\ => 
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.9\ := SmartResize(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.8\ + \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\, 64);
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_18\;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_18\ => 
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.10\ := (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.9\) < signed(SmartResize((\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num\), 64));

                        
                        
                        
                        

                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.10\) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_20\;
                        else 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_24\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_19\ => 
                        
                        
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.14\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\ + to_signed(1, 32);
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.14\;
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ = \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_19\) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_15\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_20\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.array\(to_integer(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\)).\IsNull\ := false;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.array\(to_integer(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\)).\PositBits\ := to_unsigned(0, 32);
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.11\ := SmartResize(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num3\ * to_signed(160, 32), 32);
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.12\ := to_signed(1, 32) + \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.11\;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_21\;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_21\ => 
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.13\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.12\ + \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\;
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.CellIndex\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.13\;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.ReadEnable\ <= true;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_22\;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_22\ => 
                        
                        if (\ReadsDone\ = true) then 
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.ReadEnable\ <= false;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.dataIn.1\ := \DataIn\;
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).this.parameter.Out.0\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.array\(to_integer(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\));
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).bits.parameter.Out.0\ <= ConvertStdLogicVectorToUInt32(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.dataIn.1\);
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).fromBitMask.parameter.Out.0\ <= true;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean)._Started.0\ <= true;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_23\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_23\ => 
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean)._Started.0\ = \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean)._Finished.0\) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean)._Started.0\ <= false;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.array\(to_integer(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\)) := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).this.parameter.In.0\;
                            
                            if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ = \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_23\) then 
                                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_19\;
                            end if;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_24\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.array\(to_integer(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\)).\IsNull\ := false;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.array\(to_integer(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\)).\PositBits\ := to_unsigned(0, 32);
                        
                        
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).this.parameter.Out.0\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.array\(to_integer(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\));
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).value.parameter.Out.0\ <= to_signed(0, 32);
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Started.0\ <= true;
                        \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_25\;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_25\ => 
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Started.0\ = \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Finished.0\) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Started.0\ <= false;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.array\(to_integer(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num4\)) := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).this.parameter.In.0\;
                            
                            if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ = \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_25\) then 
                                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_19\;
                            end if;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_26\ => 
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire)._Started.0\ = \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire)._Finished.0\) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire)._Started.0\ <= false;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.return.1\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).return.0\;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.array\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).posits.parameter.In.0\;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.quire\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).startingValue.parameter.In.0\;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.quire\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.return.1\;
                            
                            
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.15\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num3\ + to_signed(1, 32);
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.num3\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.binaryOperationResult.15\;
                            
                            if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ = \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_26\) then 
                                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_13\;
                            end if;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_27\ => 
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire)._Started.0\ = \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire)._Finished.0\) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire)._Started.0\ <= false;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectffd9139c321969eb0a42e1e3ae043fc0d22d96a54e32c2dc05d540c7e97af68e\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).this.parameter.In.0\;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.quire\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).q.parameter.In.0\;
                            
                            
                            
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.CellIndex\ <= to_signed(0, 32);
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.WriteEnable\ <= true;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.DataOut\ <= ConvertUInt32ToStdLogicVector(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.objectffd9139c321969eb0a42e1e3ae043fc0d22d96a54e32c2dc05d540c7e97af68e\.\PositBits\);
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_28\;
                        end if;
                        
                    when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_28\ => 
                        
                        if (\WritesDone\ = true) then 
                            
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.WriteEnable\ <= false;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State\ := \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._State_1\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::.ctor(UInt32,Boolean).0._StateMachine\: process (\Clock\) 
        Variable \Posit32::.ctor(UInt32,Boolean).0._State\: \Posit32::.ctor(UInt32,Boolean).0._States\ := \Posit32::.ctor(UInt32,Boolean).0._State_0\;
        Variable \Posit32::.ctor(UInt32,Boolean).0.this\: \Lombiq.Arithmetics.Posit32\;
        Variable \Posit32::.ctor(UInt32,Boolean).0.bits\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::.ctor(UInt32,Boolean).0.fromBitMask\: boolean := false;
        Variable \Posit32::.ctor(UInt32,Boolean).0.conditional07306ef17ce6eacdbdd521687c7db8bbabd2dc9ca02b65fce7cdbd581ebb7be6\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::.ctor(UInt32,Boolean).0._Finished\ <= false;
                \Posit32::.ctor(UInt32,Boolean).0._State\ := \Posit32::.ctor(UInt32,Boolean).0._State_0\;
                \Posit32::.ctor(UInt32,Boolean).0.bits\ := to_unsigned(0, 32);
                \Posit32::.ctor(UInt32,Boolean).0.fromBitMask\ := false;
                \Posit32::.ctor(UInt32,Boolean).0.conditional07306ef17ce6eacdbdd521687c7db8bbabd2dc9ca02b65fce7cdbd581ebb7be6\ := to_unsigned(0, 32);
            else 
                case \Posit32::.ctor(UInt32,Boolean).0._State\ is 
                    when \Posit32::.ctor(UInt32,Boolean).0._State_0\ => 
                        
                        
                        if (\Posit32::.ctor(UInt32,Boolean).0._Started\ = true) then 
                            \Posit32::.ctor(UInt32,Boolean).0._State\ := \Posit32::.ctor(UInt32,Boolean).0._State_2\;
                        end if;
                        
                    when \Posit32::.ctor(UInt32,Boolean).0._State_1\ => 
                        
                        
                        if (\Posit32::.ctor(UInt32,Boolean).0._Started\ = true) then 
                            \Posit32::.ctor(UInt32,Boolean).0._Finished\ <= true;
                        else 
                            \Posit32::.ctor(UInt32,Boolean).0._Finished\ <= false;
                            \Posit32::.ctor(UInt32,Boolean).0._State\ := \Posit32::.ctor(UInt32,Boolean).0._State_0\;
                        end if;
                        
                        \Posit32::.ctor(UInt32,Boolean).0.this.parameter.Out\ <= \Posit32::.ctor(UInt32,Boolean).0.this\;
                        
                    when \Posit32::.ctor(UInt32,Boolean).0._State_2\ => 
                        \Posit32::.ctor(UInt32,Boolean).0.this\ := \Posit32::.ctor(UInt32,Boolean).0.this.parameter.In\;
                        \Posit32::.ctor(UInt32,Boolean).0.bits\ := \Posit32::.ctor(UInt32,Boolean).0.bits.parameter.In\;
                        \Posit32::.ctor(UInt32,Boolean).0.fromBitMask\ := \Posit32::.ctor(UInt32,Boolean).0.fromBitMask.parameter.In\;
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(UInt32,Boolean).0.conditional07306ef17ce6eacdbdd521687c7db8bbabd2dc9ca02b65fce7cdbd581ebb7be6\ := \Posit32::.ctor(UInt32,Boolean).0.bits\;
                        
                        
                        
                        \Posit32::.ctor(UInt32,Boolean).0.this\.\PositBits\ := (\Posit32::.ctor(UInt32,Boolean).0.conditional07306ef17ce6eacdbdd521687c7db8bbabd2dc9ca02b65fce7cdbd581ebb7be6\);
                        \Posit32::.ctor(UInt32,Boolean).0._State\ := \Posit32::.ctor(UInt32,Boolean).0._State_1\;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::.ctor(Quire).0._StateMachine\: process (\Clock\) 
        Variable \Posit32::.ctor(Quire).0._State\: \Posit32::.ctor(Quire).0._States\ := \Posit32::.ctor(Quire).0._State_0\;
        Variable \Posit32::.ctor(Quire).0.this\: \Lombiq.Arithmetics.Posit32\;
        Variable \Posit32::.ctor(Quire).0.q\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::.ctor(Quire).0.signBit\: boolean := false;
        Variable \Posit32::.ctor(Quire).0.num\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::.ctor(Quire).0.num2\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Posit32::.ctor(Quire).0.return.0\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::.ctor(Quire).0.return.1\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.0\: boolean := false;
        Variable \Posit32::.ctor(Quire).0.return.2\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::.ctor(Quire).0.return.3\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::.ctor(Quire).0.return.4\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::.ctor(Quire).0.return.5\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.1\: boolean := false;
        Variable \Posit32::.ctor(Quire).0.return.6\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::.ctor(Quire).0.return.7\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::.ctor(Quire).0.return.8\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Posit32::.ctor(Quire).0.num3\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.3\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.4\: boolean := false;
        Variable \Posit32::.ctor(Quire).0.num4\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.5\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::.ctor(Quire).0.num5\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.6\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.7\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.8\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.9\: boolean := false;
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.10\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::.ctor(Quire).0.binaryOperationResult.11\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::.ctor(Quire).0.return.9\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::.ctor(Quire).0.return.10\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::.ctor(Quire).0.return.11\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::.ctor(Quire).0._Finished\ <= false;
                \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).right.parameter.Out.0\ <= to_signed(0, 32);
                \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ <= false;
                \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\ <= false;
                \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire)._Started.0\ <= false;
                \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).right.parameter.Out.0\ <= to_unsigned(0, 32);
                \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32)._Started.0\ <= false;
                \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\ <= to_signed(0, 32);
                \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ <= false;
                \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire)._Started.0\ <= false;
                \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).signBit.parameter.Out.0\ <= false;
                \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).regimeKValue.parameter.Out.0\ <= to_signed(0, 32);
                \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).exponentBits.parameter.Out.0\ <= to_unsigned(0, 32);
                \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).fractionBits.parameter.Out.0\ <= to_unsigned(0, 32);
                \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32)._Started.0\ <= false;
                \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_0\;
                \Posit32::.ctor(Quire).0.signBit\ := false;
                \Posit32::.ctor(Quire).0.num\ := to_signed(0, 32);
                \Posit32::.ctor(Quire).0.num2\ := to_unsigned(0, 64);
                \Posit32::.ctor(Quire).0.return.1\ := to_unsigned(0, 64);
                \Posit32::.ctor(Quire).0.binaryOperationResult.0\ := false;
                \Posit32::.ctor(Quire).0.return.5\ := to_unsigned(0, 64);
                \Posit32::.ctor(Quire).0.binaryOperationResult.1\ := false;
                \Posit32::.ctor(Quire).0.binaryOperationResult.2\ := to_signed(0, 32);
                \Posit32::.ctor(Quire).0.return.8\ := to_unsigned(0, 64);
                \Posit32::.ctor(Quire).0.num3\ := to_signed(0, 32);
                \Posit32::.ctor(Quire).0.binaryOperationResult.3\ := to_signed(0, 32);
                \Posit32::.ctor(Quire).0.binaryOperationResult.4\ := false;
                \Posit32::.ctor(Quire).0.num4\ := to_signed(0, 32);
                \Posit32::.ctor(Quire).0.binaryOperationResult.5\ := to_signed(0, 32);
                \Posit32::.ctor(Quire).0.num5\ := to_unsigned(0, 32);
                \Posit32::.ctor(Quire).0.binaryOperationResult.6\ := to_signed(0, 32);
                \Posit32::.ctor(Quire).0.binaryOperationResult.7\ := to_signed(0, 32);
                \Posit32::.ctor(Quire).0.binaryOperationResult.8\ := to_unsigned(0, 32);
                \Posit32::.ctor(Quire).0.binaryOperationResult.9\ := false;
                \Posit32::.ctor(Quire).0.binaryOperationResult.10\ := to_signed(0, 32);
                \Posit32::.ctor(Quire).0.binaryOperationResult.11\ := to_unsigned(0, 32);
                \Posit32::.ctor(Quire).0.return.10\ := to_unsigned(0, 32);
                \Posit32::.ctor(Quire).0.return.11\ := to_unsigned(0, 32);
            else 
                case \Posit32::.ctor(Quire).0._State\ is 
                    when \Posit32::.ctor(Quire).0._State_0\ => 
                        
                        
                        if (\Posit32::.ctor(Quire).0._Started\ = true) then 
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_2\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_1\ => 
                        
                        
                        if (\Posit32::.ctor(Quire).0._Started\ = true) then 
                            \Posit32::.ctor(Quire).0._Finished\ <= true;
                        else 
                            \Posit32::.ctor(Quire).0._Finished\ <= false;
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_0\;
                        end if;
                        
                        \Posit32::.ctor(Quire).0.this.parameter.Out\ <= \Posit32::.ctor(Quire).0.this\;
                        \Posit32::.ctor(Quire).0.q.parameter.Out\ <= \Posit32::.ctor(Quire).0.q\;
                        
                    when \Posit32::.ctor(Quire).0._State_2\ => 
                        \Posit32::.ctor(Quire).0.this\ := \Posit32::.ctor(Quire).0.this.parameter.In\;
                        \Posit32::.ctor(Quire).0.q\ := \Posit32::.ctor(Quire).0.q.parameter.In\;
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.this\.\PositBits\ := "10000000000000000000000000000000";
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.signBit\ := false;
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.num\ := to_signed(511, 32);
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.q\;
                        \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).right.parameter.Out.0\ <= to_signed(448, 32);
                        \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ <= true;
                        \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_3\;
                        
                    when \Posit32::.ctor(Quire).0._State_3\ => 
                        
                        if (\Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ = \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.0\ := \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).return.0\;
                            \Posit32::.ctor(Quire).0.q\ := \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.In.0\;
                            
                            \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).x.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.return.0\;
                            \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\ <= true;
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_4\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_4\ => 
                        
                        if (\Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\ = \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.1\ := \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).return.0\;
                            \Posit32::.ctor(Quire).0.return.0\ := \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).x.parameter.In.0\;
                            \Posit32::.ctor(Quire).0.num2\ := \Posit32::.ctor(Quire).0.return.1\;
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32::.ctor(Quire).0.binaryOperationResult.0\ := \Posit32::.ctor(Quire).0.num2\ >= "1000000000000000000000000000000000000000000000000000000000000000";

                            
                            
                            

                            if (\Posit32::.ctor(Quire).0.binaryOperationResult.0\) then 
                                \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_6\;
                            else 
                                
                                \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_5\;
                            end if;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_5\ => 
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.q\;
                        \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).right.parameter.Out.0\ <= to_signed(448, 32);
                        \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ <= true;
                        \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_9\;
                        
                    when \Posit32::.ctor(Quire).0._State_6\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire).q.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.q\;
                        \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire)._Started.0\ <= true;
                        \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_7\;
                        
                    when \Posit32::.ctor(Quire).0._State_7\ => 
                        
                        if (\Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire)._Started.0\ = \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.2\ := \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire).return.0\;
                            \Posit32::.ctor(Quire).0.q\ := \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire).q.parameter.In.0\;
                            \Posit32::.ctor(Quire).0.q\ := \Posit32::.ctor(Quire).0.return.2\;
                            
                            
                            
                            
                            \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).left.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.q\;
                            \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).right.parameter.Out.0\ <= to_unsigned(1, 32);
                            \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32)._Started.0\ <= true;
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_8\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_8\ => 
                        
                        if (\Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32)._Started.0\ = \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.3\ := \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).return.0\;
                            \Posit32::.ctor(Quire).0.q\ := \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).left.parameter.In.0\;
                            \Posit32::.ctor(Quire).0.q\ := \Posit32::.ctor(Quire).0.return.3\;
                            
                            
                            
                            \Posit32::.ctor(Quire).0.signBit\ := true;
                            
                            if (\Posit32::.ctor(Quire).0._State\ = \Posit32::.ctor(Quire).0._State_8\) then 
                                \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_5\;
                            end if;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_9\ => 
                        
                        if (\Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ = \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.4\ := \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).return.0\;
                            \Posit32::.ctor(Quire).0.q\ := \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.In.0\;
                            
                            \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).x.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.return.4\;
                            \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\ <= true;
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_10\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_10\ => 
                        
                        if (\Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\ = \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.5\ := \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).return.0\;
                            \Posit32::.ctor(Quire).0.return.4\ := \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).x.parameter.In.0\;
                            \Posit32::.ctor(Quire).0.num2\ := \Posit32::.ctor(Quire).0.return.5\;
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_11\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_11\ => 
                        
                        
                        
                        \Posit32::.ctor(Quire).0.binaryOperationResult.1\ := \Posit32::.ctor(Quire).0.num2\ < "1000000000000000000000000000000000000000000000000000000000000000";
                        if (\Posit32::.ctor(Quire).0.binaryOperationResult.1\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.q\;
                            \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\ <= to_signed(1, 32);
                            \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ <= true;
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_13\;
                        else 
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_12\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_12\ => 
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.binaryOperationResult.3\ := \Posit32::.ctor(Quire).0.num\ - to_signed(240, 32);
                        \Posit32::.ctor(Quire).0.num3\ := \Posit32::.ctor(Quire).0.binaryOperationResult.3\;
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.binaryOperationResult.4\ := \Posit32::.ctor(Quire).0.num\ = to_signed(0, 32);

                        
                        
                        

                        if (\Posit32::.ctor(Quire).0.binaryOperationResult.4\) then 
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_17\;
                        else 
                            
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_16\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_13\ => 
                        
                        if (\Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ = \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.6\ := \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).return.0\;
                            \Posit32::.ctor(Quire).0.q\ := \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.In.0\;
                            \Posit32::.ctor(Quire).0.q\ := \Posit32::.ctor(Quire).0.return.6\;
                            
                            
                            
                            \Posit32::.ctor(Quire).0.binaryOperationResult.2\ := \Posit32::.ctor(Quire).0.num\ - to_signed(1, 32);
                            \Posit32::.ctor(Quire).0.num\ := \Posit32::.ctor(Quire).0.binaryOperationResult.2\;
                            
                            
                            
                            
                            \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.q\;
                            \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).right.parameter.Out.0\ <= to_signed(448, 32);
                            \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ <= true;
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_14\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_14\ => 
                        
                        if (\Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ = \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.7\ := \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).return.0\;
                            \Posit32::.ctor(Quire).0.q\ := \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.In.0\;
                            
                            \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).x.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.return.7\;
                            \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\ <= true;
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_15\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_15\ => 
                        
                        if (\Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\ = \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.8\ := \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).return.0\;
                            \Posit32::.ctor(Quire).0.return.7\ := \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).x.parameter.In.0\;
                            \Posit32::.ctor(Quire).0.num2\ := \Posit32::.ctor(Quire).0.return.8\;
                            
                            if (\Posit32::.ctor(Quire).0._State\ = \Posit32::.ctor(Quire).0._State_15\) then 
                                \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_11\;
                            end if;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_16\ => 
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.binaryOperationResult.5\ := \Posit32::.ctor(Quire).0.num3\ / to_signed(4, 32);
                        \Posit32::.ctor(Quire).0.num4\ := \Posit32::.ctor(Quire).0.binaryOperationResult.5\;
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.binaryOperationResult.6\ := \Posit32::.ctor(Quire).0.num3\ / to_signed(4, 32);
                        \Posit32::.ctor(Quire).0.binaryOperationResult.7\ := SmartResize(\Posit32::.ctor(Quire).0.binaryOperationResult.6\ * to_signed(4, 32), 32);
                        \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_18\;
                        
                    when \Posit32::.ctor(Quire).0._State_17\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.this\.\PositBits\ := to_unsigned(0, 32);
                        
                        
                        
                        \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_1\;
                        
                        if (\Posit32::.ctor(Quire).0._State\ = \Posit32::.ctor(Quire).0._State_17\) then 
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_16\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_18\ => 
                        
                        \Posit32::.ctor(Quire).0.binaryOperationResult.8\ := unsigned(\Posit32::.ctor(Quire).0.num3\ - \Posit32::.ctor(Quire).0.binaryOperationResult.7\);
                        \Posit32::.ctor(Quire).0.num5\ := (\Posit32::.ctor(Quire).0.binaryOperationResult.8\);
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_19\;
                        
                    when \Posit32::.ctor(Quire).0._State_19\ => 
                        
                        \Posit32::.ctor(Quire).0.binaryOperationResult.9\ := signed(SmartResize((\Posit32::.ctor(Quire).0.num5\), 64)) < to_signed(0, 64);

                        
                        
                        

                        if (\Posit32::.ctor(Quire).0.binaryOperationResult.9\) then 
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_21\;
                        else 
                            
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_20\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_20\ => 
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.q\;
                        \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).right.parameter.Out.0\ <= to_signed(480, 32);
                        \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ <= true;
                        \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_22\;
                        
                    when \Posit32::.ctor(Quire).0._State_21\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Quire).0.binaryOperationResult.10\ := \Posit32::.ctor(Quire).0.num4\ - to_signed(1, 32);
                        \Posit32::.ctor(Quire).0.num4\ := \Posit32::.ctor(Quire).0.binaryOperationResult.10\;
                        
                        
                        
                        \Posit32::.ctor(Quire).0.binaryOperationResult.11\ := SmartResize(unsigned(signed(SmartResize((\Posit32::.ctor(Quire).0.num5\), 64)) + to_signed(4, 64)), 32);
                        \Posit32::.ctor(Quire).0.num5\ := (\Posit32::.ctor(Quire).0.binaryOperationResult.11\);
                        
                        if (\Posit32::.ctor(Quire).0._State\ = \Posit32::.ctor(Quire).0._State_21\) then 
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_20\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_22\ => 
                        
                        if (\Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ = \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.9\ := \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).return.0\;
                            \Posit32::.ctor(Quire).0.q\ := \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.In.0\;
                            
                            \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire).x.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.return.9\;
                            \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire)._Started.0\ <= true;
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_23\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_23\ => 
                        
                        if (\Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire)._Started.0\ = \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.10\ := \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire).return.0\;
                            \Posit32::.ctor(Quire).0.return.9\ := \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire).x.parameter.In.0\;
                            
                            \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).signBit.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.signBit\;
                            \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).regimeKValue.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.num4\;
                            \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).exponentBits.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.num5\;
                            \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).fractionBits.parameter.Out.0\ <= \Posit32::.ctor(Quire).0.return.10\;
                            \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32)._Started.0\ <= true;
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_24\;
                        end if;
                        
                    when \Posit32::.ctor(Quire).0._State_24\ => 
                        
                        if (\Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32)._Started.0\ = \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32)._Finished.0\) then 
                            \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32)._Started.0\ <= false;
                            \Posit32::.ctor(Quire).0.return.11\ := \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).return.0\;
                            \Posit32::.ctor(Quire).0.this\.\PositBits\ := \Posit32::.ctor(Quire).0.return.11\;
                            \Posit32::.ctor(Quire).0._State\ := \Posit32::.ctor(Quire).0._State_1\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::.ctor(UInt32).0._StateMachine\: process (\Clock\) 
        Variable \Posit32::.ctor(UInt32).0._State\: \Posit32::.ctor(UInt32).0._States\ := \Posit32::.ctor(UInt32).0._State_0\;
        Variable \Posit32::.ctor(UInt32).0.this\: \Lombiq.Arithmetics.Posit32\;
        Variable \Posit32::.ctor(UInt32).0.value\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::.ctor(UInt32).0._Finished\ <= false;
                \Posit32::.ctor(UInt32).0._State\ := \Posit32::.ctor(UInt32).0._State_0\;
                \Posit32::.ctor(UInt32).0.value\ := to_unsigned(0, 32);
            else 
                case \Posit32::.ctor(UInt32).0._State\ is 
                    when \Posit32::.ctor(UInt32).0._State_0\ => 
                        
                        
                        if (\Posit32::.ctor(UInt32).0._Started\ = true) then 
                            \Posit32::.ctor(UInt32).0._State\ := \Posit32::.ctor(UInt32).0._State_2\;
                        end if;
                        
                    when \Posit32::.ctor(UInt32).0._State_1\ => 
                        
                        
                        if (\Posit32::.ctor(UInt32).0._Started\ = true) then 
                            \Posit32::.ctor(UInt32).0._Finished\ <= true;
                        else 
                            \Posit32::.ctor(UInt32).0._Finished\ <= false;
                            \Posit32::.ctor(UInt32).0._State\ := \Posit32::.ctor(UInt32).0._State_0\;
                        end if;
                        
                        \Posit32::.ctor(UInt32).0.this.parameter.Out\ <= \Posit32::.ctor(UInt32).0.this\;
                        
                    when \Posit32::.ctor(UInt32).0._State_2\ => 
                        \Posit32::.ctor(UInt32).0.this\ := \Posit32::.ctor(UInt32).0.this.parameter.In\;
                        \Posit32::.ctor(UInt32).0.value\ := \Posit32::.ctor(UInt32).0.value.parameter.In\;
                        
                        
                        
                        \Posit32::.ctor(UInt32).0.this\.\PositBits\ := to_unsigned(0, 32);
                        \Posit32::.ctor(UInt32).0._State\ := \Posit32::.ctor(UInt32).0._State_1\;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::.ctor(Int32).0._StateMachine\: process (\Clock\) 
        Variable \Posit32::.ctor(Int32).0._State\: \Posit32::.ctor(Int32).0._States\ := \Posit32::.ctor(Int32).0._State_0\;
        Variable \Posit32::.ctor(Int32).0.this\: \Lombiq.Arithmetics.Posit32\;
        Variable \Posit32::.ctor(Int32).0.value\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::.ctor(Int32).0.conditional2430432b7cbc58715e662a8c82abb8a42239e5b92d4c7ea6c2c87a87483f3331\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::.ctor(Int32).0.object62f645adbfb4d116e9dadbde41fc03ee8eecadf80abd12f7fbc8d9dfa7162321\: \Lombiq.Arithmetics.Posit32\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::.ctor(Int32).0._Finished\ <= false;
                \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32).value.parameter.Out.0\ <= to_unsigned(0, 32);
                \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32)._Started.0\ <= false;
                \Posit32::.ctor(Int32).0._State\ := \Posit32::.ctor(Int32).0._State_0\;
                \Posit32::.ctor(Int32).0.value\ := to_signed(0, 32);
                \Posit32::.ctor(Int32).0.conditional2430432b7cbc58715e662a8c82abb8a42239e5b92d4c7ea6c2c87a87483f3331\ := to_unsigned(0, 32);
            else 
                case \Posit32::.ctor(Int32).0._State\ is 
                    when \Posit32::.ctor(Int32).0._State_0\ => 
                        
                        
                        if (\Posit32::.ctor(Int32).0._Started\ = true) then 
                            \Posit32::.ctor(Int32).0._State\ := \Posit32::.ctor(Int32).0._State_2\;
                        end if;
                        
                    when \Posit32::.ctor(Int32).0._State_1\ => 
                        
                        
                        if (\Posit32::.ctor(Int32).0._Started\ = true) then 
                            \Posit32::.ctor(Int32).0._Finished\ <= true;
                        else 
                            \Posit32::.ctor(Int32).0._Finished\ <= false;
                            \Posit32::.ctor(Int32).0._State\ := \Posit32::.ctor(Int32).0._State_0\;
                        end if;
                        
                        \Posit32::.ctor(Int32).0.this.parameter.Out\ <= \Posit32::.ctor(Int32).0.this\;
                        
                    when \Posit32::.ctor(Int32).0._State_2\ => 
                        \Posit32::.ctor(Int32).0.this\ := \Posit32::.ctor(Int32).0.this.parameter.In\;
                        \Posit32::.ctor(Int32).0.value\ := \Posit32::.ctor(Int32).0.value.parameter.In\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::.ctor(Int32).0.object62f645adbfb4d116e9dadbde41fc03ee8eecadf80abd12f7fbc8d9dfa7162321\.\IsNull\ := false;
                        \Posit32::.ctor(Int32).0.object62f645adbfb4d116e9dadbde41fc03ee8eecadf80abd12f7fbc8d9dfa7162321\.\PositBits\ := to_unsigned(0, 32);
                        
                        
                        \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32).this.parameter.Out.0\ <= \Posit32::.ctor(Int32).0.object62f645adbfb4d116e9dadbde41fc03ee8eecadf80abd12f7fbc8d9dfa7162321\;
                        \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32).value.parameter.Out.0\ <= to_unsigned(0, 32);
                        \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32)._Started.0\ <= true;
                        \Posit32::.ctor(Int32).0._State\ := \Posit32::.ctor(Int32).0._State_3\;
                        
                    when \Posit32::.ctor(Int32).0._State_3\ => 
                        
                        if (\Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32)._Started.0\ = \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32)._Finished.0\) then 
                            \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32)._Started.0\ <= false;
                            \Posit32::.ctor(Int32).0.object62f645adbfb4d116e9dadbde41fc03ee8eecadf80abd12f7fbc8d9dfa7162321\ := \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32).this.parameter.In.0\;
                            
                            
                            
                            \Posit32::.ctor(Int32).0.conditional2430432b7cbc58715e662a8c82abb8a42239e5b92d4c7ea6c2c87a87483f3331\ := to_unsigned(0, 32);
                            
                            
                            
                            \Posit32::.ctor(Int32).0.this\.\PositBits\ := to_unsigned(0, 32);
                            \Posit32::.ctor(Int32).0._State\ := \Posit32::.ctor(Int32).0._State_1\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._StateMachine\: process (\Clock\) 
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\: \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._States\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_0\;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.signBit\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.regimeKValue\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.regimeKValue_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.0\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_7433aa75d94b12689bfd37b82bd6efe2336049442f0a6f7004902fab118a3d86_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_7433aa75d94b12689bfd37b82bd6efe2336049442f0a6f7004902fab118a3d86_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b_7433aa75d94b12689bfd37b82bd6efe2336049442f0a6f7004902fab118a3d86_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.4\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.5\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.6\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.7\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.8\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.9\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.10\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.startingPosition_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.11\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.12\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.13\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.14\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.15\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.16\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.17\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.18\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.19\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.20\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.21\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.22\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.23\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional080c1e8270378fd06e215f3c8f2add99c4865c1fbe8dd647a36c0c7e2edafab9\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.24\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.25\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.26\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.27\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.28\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional8ec324176b3f3fcd58fd5cfa6806fcab9222414090d26d94c66a65f1e77ad791\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.29\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.30\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.31\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.32\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.33\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.34\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalc44e6e18dba54d497a9ebfd5cd45c62d920ed273ec5aec35f89d9d27a8e797d3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_29d01fc597480c9a8978df84b3fa377f862967419a63789112fc92c8bcb8358e\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_29d01fc597480c9a8978df84b3fa377f862967419a63789112fc92c8bcb8358e\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.35\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalfaf425f73af9abdd07507acc85c797211aab0cbc36083f9065056c957f27c6b3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.36\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.37\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.38\: signed(63 downto 0) := to_signed(0, 64);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.39\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalb43e86d5d828dd5119f9f88af0ba7c790398b5cca8ee395bf1a45e5780b616e0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_c365944f32d1bd43cad8b7e282704038c75bff2f7f5617940490de000fbf3f9f\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_c365944f32d1bd43cad8b7e282704038c75bff2f7f5617940490de000fbf3f9f\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.40\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num3\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_3938d622f1c7059e43ce720914f8dac78e0c43b14e9f57ead44226443ac08a49\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_3938d622f1c7059e43ce720914f8dac78e0c43b14e9f57ead44226443ac08a49\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b_3938d622f1c7059e43ce720914f8dac78e0c43b14e9f57ead44226443ac08a49\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.41\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.42\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.43\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.44\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_1f023f1605903ad9d771877041978dfe685eea174a0d8f4cd7264316130e8abc\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.index_1f023f1605903ad9d771877041978dfe685eea174a0d8f4cd7264316130e8abc\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_1f023f1605903ad9d771877041978dfe685eea174a0d8f4cd7264316130e8abc\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.45\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.4\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.46\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num4\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.47\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.48\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalbf654792f1ef201c91607ce88a255151da71234b0142c97b5e2a3594fec8b3f2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.49\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.50\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.5\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.51\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.52\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.53\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional0557e32b11ba8656de63af77389f74397db38458b6838b7ec71d9300b43b97b3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.54\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.55\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.56\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.6\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.57\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.58\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.59\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.60\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional18df916b486c957f6d73b71f963f462865051a4dad21055f9f7bb67a1b272e87\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.61\: boolean := false;
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.62\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.63\: signed(63 downto 0) := to_signed(0, 64);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.64\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionala777843480080cfd7ce563a33d79f12dd3aff5a7f1e7ee2bc6ae68dce3ba9f02\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_d5e78a1cc4c5ce9ecd46e134cd314afbdaeeeb0c6ac7678364f0a765152de487\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_d5e78a1cc4c5ce9ecd46e134cd314afbdaeeeb0c6ac7678364f0a765152de487\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.7\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.65\: unsigned(31 downto 0) := to_unsigned(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._Finished\ <= false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return\ <= to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_0\;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.signBit\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.regimeKValue\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.regimeKValue_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.0\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.1\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.2\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.3\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_7433aa75d94b12689bfd37b82bd6efe2336049442f0a6f7004902fab118a3d86_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_7433aa75d94b12689bfd37b82bd6efe2336049442f0a6f7004902fab118a3d86_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\ := to_unsigned(0, 8);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b_7433aa75d94b12689bfd37b82bd6efe2336049442f0a6f7004902fab118a3d86_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\ := to_unsigned(0, 8);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.4\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.5\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.6\ := to_unsigned(0, 8);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.7\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.8\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.9\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.0\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.10\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b\ := to_unsigned(0, 8);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.startingPosition_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\ := to_unsigned(0, 8);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\ := to_unsigned(0, 8);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\ := to_unsigned(0, 8);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.11\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.12\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.13\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.14\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.15\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.16\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.17\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.18\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.19\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.20\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.21\ := to_unsigned(0, 8);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.22\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.23\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional080c1e8270378fd06e215f3c8f2add99c4865c1fbe8dd647a36c0c7e2edafab9\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.24\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.25\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.1\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.26\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.27\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.28\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional8ec324176b3f3fcd58fd5cfa6806fcab9222414090d26d94c66a65f1e77ad791\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.29\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.30\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.31\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.32\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.33\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.34\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalc44e6e18dba54d497a9ebfd5cd45c62d920ed273ec5aec35f89d9d27a8e797d3\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_29d01fc597480c9a8978df84b3fa377f862967419a63789112fc92c8bcb8358e\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_29d01fc597480c9a8978df84b3fa377f862967419a63789112fc92c8bcb8358e\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.2\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.35\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalfaf425f73af9abdd07507acc85c797211aab0cbc36083f9065056c957f27c6b3\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.36\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.37\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.38\ := to_signed(0, 64);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.39\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalb43e86d5d828dd5119f9f88af0ba7c790398b5cca8ee395bf1a45e5780b616e0\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_c365944f32d1bd43cad8b7e282704038c75bff2f7f5617940490de000fbf3f9f\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_c365944f32d1bd43cad8b7e282704038c75bff2f7f5617940490de000fbf3f9f\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.3\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.40\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num3\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_3938d622f1c7059e43ce720914f8dac78e0c43b14e9f57ead44226443ac08a49\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_3938d622f1c7059e43ce720914f8dac78e0c43b14e9f57ead44226443ac08a49\ := to_unsigned(0, 8);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b_3938d622f1c7059e43ce720914f8dac78e0c43b14e9f57ead44226443ac08a49\ := to_unsigned(0, 8);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.41\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.42\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.43\ := to_unsigned(0, 8);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.44\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_1f023f1605903ad9d771877041978dfe685eea174a0d8f4cd7264316130e8abc\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.index_1f023f1605903ad9d771877041978dfe685eea174a0d8f4cd7264316130e8abc\ := to_unsigned(0, 16);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_1f023f1605903ad9d771877041978dfe685eea174a0d8f4cd7264316130e8abc\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.45\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.4\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.46\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num4\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.47\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.48\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalbf654792f1ef201c91607ce88a255151da71234b0142c97b5e2a3594fec8b3f2\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.49\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.50\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.5\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.51\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.52\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.53\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional0557e32b11ba8656de63af77389f74397db38458b6838b7ec71d9300b43b97b3\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.54\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.55\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.56\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.6\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.57\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.58\ := to_signed(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.59\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.60\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional18df916b486c957f6d73b71f963f462865051a4dad21055f9f7bb67a1b272e87\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.61\ := false;
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.62\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.63\ := to_signed(0, 64);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.64\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionala777843480080cfd7ce563a33d79f12dd3aff5a7f1e7ee2bc6ae68dce3ba9f02\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_d5e78a1cc4c5ce9ecd46e134cd314afbdaeeeb0c6ac7678364f0a765152de487\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_d5e78a1cc4c5ce9ecd46e134cd314afbdaeeeb0c6ac7678364f0a765152de487\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.7\ := to_unsigned(0, 32);
                \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.65\ := to_unsigned(0, 32);
            else 
                case \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ is 
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_0\ => 
                        
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._Started\ = true) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_2\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_1\ => 
                        
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._Started\ = true) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._Finished\ <= true;
                        else 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._Finished\ <= false;
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_0\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_2\ => 
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.signBit\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.signBit.parameter.In\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.regimeKValue\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.regimeKValue.parameter.In\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits.parameter.In\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits.parameter.In\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.regimeKValue_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.regimeKValue\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.0\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.regimeKValue_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\ > to_signed(0, 32);

                        
                        
                        

                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.0\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_5\;
                        else 
                            
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_4\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_3\ => 
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\;
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.startingPosition_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\ := SmartResize(unsigned(to_signed(31, 32)), 8);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\ := SmartResize(unsigned(to_signed(1, 32)), 8);
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.11\ := to_signed(32, 32) - signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.startingPosition_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\), 32));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.12\ := shift_left(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\, to_integer(unsigned(SmartResize(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.11\, 5))));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.12\;
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_12\;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_4\ => 
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.0\ := -\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.regimeKValue_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.10\ := shift_right(to_unsigned(1073741824, 32), to_integer(unsigned(SmartResize(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.0\, 5) and "11111")));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.10\;
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_3\;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_5\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.1\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.regimeKValue_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\ + to_signed(1, 32);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.2\ := shift_left(to_signed(1, 32), to_integer(unsigned(SmartResize(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.1\, 5))));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_6\;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_6\ => 
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.3\ := unsigned((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.2\) - to_signed(1, 32));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.3\);
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_7433aa75d94b12689bfd37b82bd6efe2336049442f0a6f7004902fab118a3d86_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b_7433aa75d94b12689bfd37b82bd6efe2336049442f0a6f7004902fab118a3d86_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\ := SmartResize(unsigned(to_signed(0, 32)), 8);
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_7\;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_7\ => 
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.4\ := signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_7433aa75d94b12689bfd37b82bd6efe2336049442f0a6f7004902fab118a3d86_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\), 64)) /= to_signed(0, 64);
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.4\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.5\ := shift_right(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_7433aa75d94b12689bfd37b82bd6efe2336049442f0a6f7004902fab118a3d86_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\, to_integer(unsigned(SmartResize(to_signed(1, 32), 5) and "11111")));
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_7433aa75d94b12689bfd37b82bd6efe2336049442f0a6f7004902fab118a3d86_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.5\;
                            
                            
                            
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_9\;
                        else 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_8\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_8\ => 
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_7433aa75d94b12689bfd37b82bd6efe2336049442f0a6f7004902fab118a3d86_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b_7433aa75d94b12689bfd37b82bd6efe2336049442f0a6f7004902fab118a3d86_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\;
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.7\ := to_signed(32, 32) - signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_7433aa75d94b12689bfd37b82bd6efe2336049442f0a6f7004902fab118a3d86_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\), 32));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.8\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.7\ - to_signed(1, 32);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_10\;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_9\ => 
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.6\ := SmartResize(unsigned(signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b_7433aa75d94b12689bfd37b82bd6efe2336049442f0a6f7004902fab118a3d86_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\), 32)) + to_signed(1, 32)), 8);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b_7433aa75d94b12689bfd37b82bd6efe2336049442f0a6f7004902fab118a3d86_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.6\);
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_9\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_7\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_10\ => 
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.9\ := shift_left(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\, to_integer(unsigned(SmartResize(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.8\, 5))));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_877cc8a4458b184cbefcdd364edb21dd8da2ca93f5d0907ebe0e479c950d39da\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.9\;
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_3\;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_11\ => 
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_11\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_4\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_12\ => 
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.13\ := shift_right(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\, to_integer(unsigned(SmartResize(to_signed(31, 32), 5) and "11111")));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.14\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.13\) and to_unsigned(1, 32);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.14\;
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.15\ := shift_left(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\, to_integer(unsigned(SmartResize(to_signed(1, 32), 5))));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.15\;
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\ := to_signed(0, 32);
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_13\;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_13\ => 
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.16\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\) < signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.startingPosition_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\), 32));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.17\ := shift_right(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\, to_integer(unsigned(SmartResize(to_signed(31, 32), 5) and "11111")));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_15\;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_14\ => 
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\;
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\;
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.23\ := to_signed(28, 32) - signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b\), 32));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.23\);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.24\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2\ >= to_signed(0, 32);

                        
                        
                        
                        

                        if ((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.24\)) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_18\;
                        else 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_19\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_15\ => 
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.18\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.17\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.19\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.16\ and \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.18\;
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.19\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.20\ := shift_left(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\, to_integer(unsigned(SmartResize(to_signed(1, 32), 5))));
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.20\;
                            
                            
                            
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_16\;
                        else 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_14\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_16\ => 
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.21\ := SmartResize(unsigned(signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\), 32)) + to_signed(1, 32)), 8);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.21\);
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.22\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\ + to_signed(1, 32);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2_1a2fe290ae47b1ef7ded540ce3403c2e5603c310223a0b07c1ac70a272d6301b\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.22\;
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_16\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_13\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_17\ => 
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.27\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\ + (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional080c1e8270378fd06e215f3c8f2add99c4865c1fbe8dd647a36c0c7e2edafab9\);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.27\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.28\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2\ < to_signed(0, 32);

                        
                        
                        

                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.28\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_21\;
                        else 
                            
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_20\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_18\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.25\ := shift_left(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits\, to_integer(unsigned(SmartResize(unsigned(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2\), 5))));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional080c1e8270378fd06e215f3c8f2add99c4865c1fbe8dd647a36c0c7e2edafab9\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.25\);
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_18\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_17\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_19\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.1\ := -\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.26\ := shift_right(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits\, to_integer(unsigned(SmartResize(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.1\, 5) and "11111")));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional080c1e8270378fd06e215f3c8f2add99c4865c1fbe8dd647a36c0c7e2edafab9\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.26\);
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_19\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_17\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_20\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_3938d622f1c7059e43ce720914f8dac78e0c43b14e9f57ead44226443ac08a49\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b_3938d622f1c7059e43ce720914f8dac78e0c43b14e9f57ead44226443ac08a49\ := SmartResize(unsigned(to_signed(0, 32)), 8);
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_37\;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_21\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.29\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2\ > to_signed(28, 32);

                        
                        
                        
                        

                        if ((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.29\)) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_23\;
                        else 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_25\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_22\ => 
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional8ec324176b3f3fcd58fd5cfa6806fcab9222414090d26d94c66a65f1e77ad791\);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.34\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits\ < "10000000000000000000000000000000";

                        
                        
                        

                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.34\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_27\;
                        else 
                            
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_26\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_23\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.30\ := to_signed(32, 32) + \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_24\;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_24\ => 
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.31\ := shift_right(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits\, to_integer(unsigned(SmartResize(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.30\, 5) and "11111")));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional8ec324176b3f3fcd58fd5cfa6806fcab9222414090d26d94c66a65f1e77ad791\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.31\);
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_24\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_22\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_25\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.32\ := to_signed(32, 32) + \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num2\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.33\ := shift_left(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits\, to_integer(unsigned(SmartResize(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.32\, 5))));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional8ec324176b3f3fcd58fd5cfa6806fcab9222414090d26d94c66a65f1e77ad791\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.33\);
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_25\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_22\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_26\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.36\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits\ /= "10000000000000000000000000000000";

                        
                        
                        
                        

                        if ((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.36\)) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_32\;
                        else 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_33\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_27\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        

                        
                        
                        
                        

                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.signBit\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_29\;
                        else 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_30\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_28\ => 
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalc44e6e18dba54d497a9ebfd5cd45c62d920ed273ec5aec35f89d9d27a8e797d3\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_1\;
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_28\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_26\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_29\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_29d01fc597480c9a8978df84b3fa377f862967419a63789112fc92c8bcb8358e\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\;
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.2\ := not(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_29d01fc597480c9a8978df84b3fa377f862967419a63789112fc92c8bcb8358e\);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.35\ := SmartResize(unsigned(signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.2\), 64)) + to_signed(1, 64)), 32);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_29d01fc597480c9a8978df84b3fa377f862967419a63789112fc92c8bcb8358e\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.35\);
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalc44e6e18dba54d497a9ebfd5cd45c62d920ed273ec5aec35f89d9d27a8e797d3\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_29d01fc597480c9a8978df84b3fa377f862967419a63789112fc92c8bcb8358e\;
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_29\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_28\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_30\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalc44e6e18dba54d497a9ebfd5cd45c62d920ed273ec5aec35f89d9d27a8e797d3\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\;
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_30\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_28\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_31\ => 
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalfaf425f73af9abdd07507acc85c797211aab0cbc36083f9065056c957f27c6b3\);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        

                        
                        
                        
                        

                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.signBit\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_35\;
                        else 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_36\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_32\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.37\ := SmartResize(unsigned(signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\), 64)) + to_signed(1, 64)), 32);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalfaf425f73af9abdd07507acc85c797211aab0cbc36083f9065056c957f27c6b3\ := ((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.37\));
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_32\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_31\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_33\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.38\ := signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\), 64)) and to_signed(1, 64);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.39\ := SmartResize(unsigned(signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\), 64)) + (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.38\)), 32);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalfaf425f73af9abdd07507acc85c797211aab0cbc36083f9065056c957f27c6b3\ := ((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.39\));
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_33\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_31\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_34\ => 
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalb43e86d5d828dd5119f9f88af0ba7c790398b5cca8ee395bf1a45e5780b616e0\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_1\;
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_34\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_20\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_35\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_c365944f32d1bd43cad8b7e282704038c75bff2f7f5617940490de000fbf3f9f\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\;
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.3\ := not(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_c365944f32d1bd43cad8b7e282704038c75bff2f7f5617940490de000fbf3f9f\);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.40\ := SmartResize(unsigned(signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.3\), 64)) + to_signed(1, 64)), 32);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_c365944f32d1bd43cad8b7e282704038c75bff2f7f5617940490de000fbf3f9f\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.40\);
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalb43e86d5d828dd5119f9f88af0ba7c790398b5cca8ee395bf1a45e5780b616e0\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_c365944f32d1bd43cad8b7e282704038c75bff2f7f5617940490de000fbf3f9f\;
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_35\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_34\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_36\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalb43e86d5d828dd5119f9f88af0ba7c790398b5cca8ee395bf1a45e5780b616e0\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\;
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_36\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_34\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_37\ => 
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.41\ := signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_3938d622f1c7059e43ce720914f8dac78e0c43b14e9f57ead44226443ac08a49\), 64)) /= to_signed(0, 64);
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.41\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.42\ := shift_right(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_3938d622f1c7059e43ce720914f8dac78e0c43b14e9f57ead44226443ac08a49\, to_integer(unsigned(SmartResize(to_signed(1, 32), 5) and "11111")));
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_3938d622f1c7059e43ce720914f8dac78e0c43b14e9f57ead44226443ac08a49\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.42\;
                            
                            
                            
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_39\;
                        else 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_38\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_38\ => 
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_3938d622f1c7059e43ce720914f8dac78e0c43b14e9f57ead44226443ac08a49\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b_3938d622f1c7059e43ce720914f8dac78e0c43b14e9f57ead44226443ac08a49\;
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.44\ := signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_3938d622f1c7059e43ce720914f8dac78e0c43b14e9f57ead44226443ac08a49\), 32)) - to_signed(1, 32);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num3\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.44\);
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_1f023f1605903ad9d771877041978dfe685eea174a0d8f4cd7264316130e8abc\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\;
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.index_1f023f1605903ad9d771877041978dfe685eea174a0d8f4cd7264316130e8abc\ := SmartResize(unsigned(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num3\), 16);
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.45\ := shift_left(to_signed(1, 32), to_integer(unsigned(SmartResize(signed(SmartResize(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.index_1f023f1605903ad9d771877041978dfe685eea174a0d8f4cd7264316130e8abc\, 32)), 5))));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.4\ := not((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.45\));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_40\;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_39\ => 
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.43\ := SmartResize(unsigned(signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b_3938d622f1c7059e43ce720914f8dac78e0c43b14e9f57ead44226443ac08a49\), 32)) + to_signed(1, 32)), 8);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b_3938d622f1c7059e43ce720914f8dac78e0c43b14e9f57ead44226443ac08a49\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.43\);
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_39\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_37\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_40\ => 
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.46\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_1f023f1605903ad9d771877041978dfe685eea174a0d8f4cd7264316130e8abc\ and unsigned((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.4\));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_1f023f1605903ad9d771877041978dfe685eea174a0d8f4cd7264316130e8abc\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.46\;
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_1f023f1605903ad9d771877041978dfe685eea174a0d8f4cd7264316130e8abc\;
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.47\ := to_signed(28, 32) - \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num3\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.48\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.47\) - signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.b\), 32));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num4\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.48\);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_41\;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_41\ => 
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.49\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num4\ >= to_signed(0, 32);

                        
                        
                        
                        

                        if ((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.49\)) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_43\;
                        else 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_44\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_42\ => 
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.52\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\ + (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalbf654792f1ef201c91607ce88a255151da71234b0142c97b5e2a3594fec8b3f2\);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.52\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.53\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num4\ < to_signed(0, 32);

                        
                        
                        

                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.53\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_46\;
                        else 
                            
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_45\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_43\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.50\ := shift_left(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\, to_integer(unsigned(SmartResize(unsigned(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num4\), 5))));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalbf654792f1ef201c91607ce88a255151da71234b0142c97b5e2a3594fec8b3f2\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.50\);
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_43\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_42\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_44\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.5\ := -\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num4\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.51\ := shift_right(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\, to_integer(unsigned(SmartResize(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.5\, 5) and "11111")));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionalbf654792f1ef201c91607ce88a255151da71234b0142c97b5e2a3594fec8b3f2\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.51\);
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_44\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_42\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_45\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        

                        
                        
                        
                        

                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.signBit\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_57\;
                        else 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_58\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_46\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.54\ := to_signed(32, 32) + \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num4\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.55\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.54\ < to_signed(0, 32);

                        
                        
                        
                        

                        if ((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.55\)) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_48\;
                        else 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_50\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_47\ => 
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional0557e32b11ba8656de63af77389f74397db38458b6838b7ec71d9300b43b97b3\);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.60\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\ >= "10000000000000000000000000000000";

                        
                        
                        

                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.60\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_52\;
                        else 
                            
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_51\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_48\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.56\ := to_signed(32, 32) - \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num4\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.6\ := -(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.56\);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_49\;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_49\ => 
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.57\ := shift_right(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\, to_integer(unsigned(SmartResize(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.6\, 5) and "11111")));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional0557e32b11ba8656de63af77389f74397db38458b6838b7ec71d9300b43b97b3\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.57\);
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_49\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_47\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_50\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.58\ := to_signed(32, 32) + \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num4\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.59\ := shift_left(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\, to_integer(unsigned(SmartResize(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.58\, 5))));
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional0557e32b11ba8656de63af77389f74397db38458b6838b7ec71d9300b43b97b3\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.59\);
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_50\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_47\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_51\ => 
                        
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_51\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_45\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_52\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.61\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits\ /= "10000000000000000000000000000000";

                        
                        
                        
                        

                        if ((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.61\)) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_54\;
                        else 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_55\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_53\ => 
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional18df916b486c957f6d73b71f963f462865051a4dad21055f9f7bb67a1b272e87\);
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_53\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_51\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_54\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.62\ := SmartResize(unsigned(signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\), 64)) + to_signed(1, 64)), 32);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional18df916b486c957f6d73b71f963f462865051a4dad21055f9f7bb67a1b272e87\ := ((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.62\));
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_54\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_53\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_55\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.63\ := signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\), 64)) and to_signed(1, 64);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.64\ := SmartResize(unsigned(signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\), 64)) + (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.63\)), 32);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditional18df916b486c957f6d73b71f963f462865051a4dad21055f9f7bb67a1b272e87\ := ((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.64\));
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_55\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_53\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_56\ => 
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionala777843480080cfd7ce563a33d79f12dd3aff5a7f1e7ee2bc6ae68dce3ba9f02\;
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_1\;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_57\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_d5e78a1cc4c5ce9ecd46e134cd314afbdaeeeb0c6ac7678364f0a765152de487\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\;
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.7\ := not(\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.bits_d5e78a1cc4c5ce9ecd46e134cd314afbdaeeeb0c6ac7678364f0a765152de487\);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.65\ := SmartResize(unsigned(signed(SmartResize((\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.unaryOperationResult.7\), 64)) + to_signed(1, 64)), 32);
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_d5e78a1cc4c5ce9ecd46e134cd314afbdaeeeb0c6ac7678364f0a765152de487\ := (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.binaryOperationResult.65\);
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionala777843480080cfd7ce563a33d79f12dd3aff5a7f1e7ee2bc6ae68dce3ba9f02\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return_d5e78a1cc4c5ce9ecd46e134cd314afbdaeeeb0c6ac7678364f0a765152de487\;
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_57\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_56\;
                        end if;
                        
                    when \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_58\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.conditionala777843480080cfd7ce563a33d79f12dd3aff5a7f1e7ee2bc6ae68dce3ba9f02\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.num\;
                        
                        if (\Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ = \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_58\) then 
                            \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State\ := \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._State_56\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Posit32::FusedSum(Posit32[],Quire).0._StateMachine\: process (\Clock\) 
        Variable \Posit32::FusedSum(Posit32[],Quire).0._State\: \Posit32::FusedSum(Posit32[],Quire).0._States\ := \Posit32::FusedSum(Posit32[],Quire).0._State_0\;
        Variable \Posit32::FusedSum(Posit32[],Quire).0.posits\: \Lombiq.Arithmetics.Posit32_Array\(0 to 159);
        Variable \Posit32::FusedSum(Posit32[],Quire).0.startingValue\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::FusedSum(Posit32[],Quire).0.quire\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::FusedSum(Posit32[],Quire).0.objectcca0dec009ae8ed2326a07122a465f3ec1a2db6344ea5f25f4320f84fc89c011\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::FusedSum(Posit32[],Quire).0.return.0\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::FusedSum(Posit32[],Quire).0.return.1\: boolean := false;
        Variable \Posit32::FusedSum(Posit32[],Quire).0.num\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Posit32::FusedSum(Posit32[],Quire).0.binaryOperationResult.0\: boolean := false;
        Variable \Posit32::FusedSum(Posit32[],Quire).0.this_5a35665db2c694b12f0378313997a8c2bfbceb9e55e0f30abbc5b3e06d2ec2d4\: \Lombiq.Arithmetics.Posit32\;
        Variable \Posit32::FusedSum(Posit32[],Quire).0.return_5a35665db2c694b12f0378313997a8c2bfbceb9e55e0f30abbc5b3e06d2ec2d4\: boolean := false;
        Variable \Posit32::FusedSum(Posit32[],Quire).0.binaryOperationResult.1\: boolean := false;
        Variable \Posit32::FusedSum(Posit32[],Quire).0.return.2\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::FusedSum(Posit32[],Quire).0.return.3\: \Lombiq.Arithmetics.Quire\;
        Variable \Posit32::FusedSum(Posit32[],Quire).0.binaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Posit32::FusedSum(Posit32[],Quire).0._Finished\ <= false;
                \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).firstSegment.parameter.Out.0\ <= to_unsigned(0, 32);
                \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Started.0\ <= false;
                \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\ <= to_signed(0, 32);
                \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ <= false;
                \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire)._Started.0\ <= false;
                \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Started.0\ <= false;
                \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\ <= false;
                \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_0\;
                \Posit32::FusedSum(Posit32[],Quire).0.return.1\ := false;
                \Posit32::FusedSum(Posit32[],Quire).0.num\ := to_signed(0, 32);
                \Posit32::FusedSum(Posit32[],Quire).0.binaryOperationResult.0\ := false;
                \Posit32::FusedSum(Posit32[],Quire).0.return_5a35665db2c694b12f0378313997a8c2bfbceb9e55e0f30abbc5b3e06d2ec2d4\ := false;
                \Posit32::FusedSum(Posit32[],Quire).0.binaryOperationResult.1\ := false;
                \Posit32::FusedSum(Posit32[],Quire).0.binaryOperationResult.2\ := to_signed(0, 32);
            else 
                case \Posit32::FusedSum(Posit32[],Quire).0._State\ is 
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_0\ => 
                        
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0._Started\ = true) then 
                            \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_2\;
                        end if;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_1\ => 
                        
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0._Started\ = true) then 
                            \Posit32::FusedSum(Posit32[],Quire).0._Finished\ <= true;
                        else 
                            \Posit32::FusedSum(Posit32[],Quire).0._Finished\ <= false;
                            \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_0\;
                        end if;
                        
                        \Posit32::FusedSum(Posit32[],Quire).0.posits.parameter.Out\ <= \Posit32::FusedSum(Posit32[],Quire).0.posits\;
                        \Posit32::FusedSum(Posit32[],Quire).0.startingValue.parameter.Out\ <= \Posit32::FusedSum(Posit32[],Quire).0.startingValue\;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_2\ => 
                        \Posit32::FusedSum(Posit32[],Quire).0.posits\ := \Posit32::FusedSum(Posit32[],Quire).0.posits.parameter.In\;
                        \Posit32::FusedSum(Posit32[],Quire).0.startingValue\ := \Posit32::FusedSum(Posit32[],Quire).0.startingValue.parameter.In\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::FusedSum(Posit32[],Quire).0.objectcca0dec009ae8ed2326a07122a465f3ec1a2db6344ea5f25f4320f84fc89c011\.\IsNull\ := false;
                        \Posit32::FusedSum(Posit32[],Quire).0.objectcca0dec009ae8ed2326a07122a465f3ec1a2db6344ea5f25f4320f84fc89c011\.\Size\ := to_unsigned(0, 16);
                        \Posit32::FusedSum(Posit32[],Quire).0.objectcca0dec009ae8ed2326a07122a465f3ec1a2db6344ea5f25f4320f84fc89c011\.\SegmentCount\ := to_unsigned(0, 16);
                        \Posit32::FusedSum(Posit32[],Quire).0.objectcca0dec009ae8ed2326a07122a465f3ec1a2db6344ea5f25f4320f84fc89c011\.\Segments\ := (others => to_unsigned(0, 64));
                        
                        
                        \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).this.parameter.Out.0\ <= \Posit32::FusedSum(Posit32[],Quire).0.objectcca0dec009ae8ed2326a07122a465f3ec1a2db6344ea5f25f4320f84fc89c011\;
                        \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).firstSegment.parameter.Out.0\ <= to_unsigned(1, 32);
                        \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).size.parameter.Out.0\ <= SmartResize(unsigned(to_signed(512, 32)), 16);
                        \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Started.0\ <= true;
                        \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_3\;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_3\ => 
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Started.0\ = \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Finished.0\) then 
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Started.0\ <= false;
                            \Posit32::FusedSum(Posit32[],Quire).0.objectcca0dec009ae8ed2326a07122a465f3ec1a2db6344ea5f25f4320f84fc89c011\ := \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).this.parameter.In.0\;
                            
                            
                            
                            
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.Out.0\ <= \Posit32::FusedSum(Posit32[],Quire).0.objectcca0dec009ae8ed2326a07122a465f3ec1a2db6344ea5f25f4320f84fc89c011\;
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\ <= to_signed(511, 32);
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ <= true;
                            \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_4\;
                        end if;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_4\ => 
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ = \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\) then 
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ <= false;
                            \Posit32::FusedSum(Posit32[],Quire).0.return.0\ := \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).return.0\;
                            \Posit32::FusedSum(Posit32[],Quire).0.objectcca0dec009ae8ed2326a07122a465f3ec1a2db6344ea5f25f4320f84fc89c011\ := \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.In.0\;
                            \Posit32::FusedSum(Posit32[],Quire).0.quire\ := \Posit32::FusedSum(Posit32[],Quire).0.return.0\;
                            
                            
                            
                            
                            
                            
                            \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).left.parameter.Out.0\ <= \Posit32::FusedSum(Posit32[],Quire).0.startingValue\;
                            \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).right.parameter.Out.0\ <= \Posit32::FusedSum(Posit32[],Quire).0.quire\;
                            \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire)._Started.0\ <= true;
                            \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_5\;
                        end if;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_5\ => 
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire)._Started.0\ = \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire)._Finished.0\) then 
                            \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire)._Started.0\ <= false;
                            \Posit32::FusedSum(Posit32[],Quire).0.return.1\ := \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).return.0\;
                            \Posit32::FusedSum(Posit32[],Quire).0.startingValue\ := \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).left.parameter.In.0\;
                            \Posit32::FusedSum(Posit32[],Quire).0.quire\ := \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).right.parameter.In.0\;

                            
                            
                            

                            if (\Posit32::FusedSum(Posit32[],Quire).0.return.1\) then 
                                \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_7\;
                            else 
                                
                                \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_6\;
                            end if;
                        end if;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_6\ => 
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::FusedSum(Posit32[],Quire).0.num\ := to_signed(0, 32);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_8\;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_7\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::FusedSum(Posit32[],Quire).0.return\ <= \Posit32::FusedSum(Posit32[],Quire).0.quire\;
                        \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_1\;
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0._State\ = \Posit32::FusedSum(Posit32[],Quire).0._State_7\) then 
                            \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_6\;
                        end if;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_8\ => 
                        
                        
                        \Posit32::FusedSum(Posit32[],Quire).0.binaryOperationResult.0\ := \Posit32::FusedSum(Posit32[],Quire).0.num\ < to_signed(160, 32);
                        if (\Posit32::FusedSum(Posit32[],Quire).0.binaryOperationResult.0\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32::FusedSum(Posit32[],Quire).0.this_5a35665db2c694b12f0378313997a8c2bfbceb9e55e0f30abbc5b3e06d2ec2d4\ := \Posit32::FusedSum(Posit32[],Quire).0.posits\(to_integer(\Posit32::FusedSum(Posit32[],Quire).0.num\));
                            
                            
                            
                            
                            
                            
                            
                            
                            \Posit32::FusedSum(Posit32[],Quire).0.binaryOperationResult.1\ := \Posit32::FusedSum(Posit32[],Quire).0.this_5a35665db2c694b12f0378313997a8c2bfbceb9e55e0f30abbc5b3e06d2ec2d4\.\PositBits\ = "10000000000000000000000000000000";
                            \Posit32::FusedSum(Posit32[],Quire).0.return_5a35665db2c694b12f0378313997a8c2bfbceb9e55e0f30abbc5b3e06d2ec2d4\ := \Posit32::FusedSum(Posit32[],Quire).0.binaryOperationResult.1\;
                            
                            
                            
                            
                            

                            
                            
                            

                            if (\Posit32::FusedSum(Posit32[],Quire).0.return_5a35665db2c694b12f0378313997a8c2bfbceb9e55e0f30abbc5b3e06d2ec2d4\) then 
                                \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_11\;
                            else 
                                
                                \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_10\;
                            end if;
                        else 
                            \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_9\;
                        end if;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_9\ => 
                        
                        
                        
                        
                        \Posit32::FusedSum(Posit32[],Quire).0.return\ <= \Posit32::FusedSum(Posit32[],Quire).0.startingValue\;
                        \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_1\;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_10\ => 
                        
                        
                        
                        
                        
                        \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32).x.parameter.Out.0\ <= \Posit32::FusedSum(Posit32[],Quire).0.posits\(to_integer(\Posit32::FusedSum(Posit32[],Quire).0.num\));
                        \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Started.0\ <= true;
                        \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_12\;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_11\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Posit32::FusedSum(Posit32[],Quire).0.return\ <= \Posit32::FusedSum(Posit32[],Quire).0.quire\;
                        \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_1\;
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0._State\ = \Posit32::FusedSum(Posit32[],Quire).0._State_11\) then 
                            \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_10\;
                        end if;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_12\ => 
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Started.0\ = \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\) then 
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Started.0\ <= false;
                            \Posit32::FusedSum(Posit32[],Quire).0.return.2\ := \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32).return.0\;
                            
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.Out.0\ <= \Posit32::FusedSum(Posit32[],Quire).0.startingValue\;
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.Out.0\ <= \Posit32::FusedSum(Posit32[],Quire).0.return.2\;
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\ <= true;
                            \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_13\;
                        end if;
                        
                    when \Posit32::FusedSum(Posit32[],Quire).0._State_13\ => 
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\ = \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\) then 
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\ <= false;
                            \Posit32::FusedSum(Posit32[],Quire).0.return.3\ := \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).return.0\;
                            \Posit32::FusedSum(Posit32[],Quire).0.startingValue\ := \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.In.0\;
                            \Posit32::FusedSum(Posit32[],Quire).0.return.2\ := \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.In.0\;
                            \Posit32::FusedSum(Posit32[],Quire).0.startingValue\ := \Posit32::FusedSum(Posit32[],Quire).0.return.3\;
                            
                            
                            
                            \Posit32::FusedSum(Posit32[],Quire).0.binaryOperationResult.2\ := \Posit32::FusedSum(Posit32[],Quire).0.num\ + to_signed(1, 32);
                            \Posit32::FusedSum(Posit32[],Quire).0.num\ := \Posit32::FusedSum(Posit32[],Quire).0.binaryOperationResult.2\;
                            
                            if (\Posit32::FusedSum(Posit32[],Quire).0._State\ = \Posit32::FusedSum(Posit32[],Quire).0._State_13\) then 
                                \Posit32::FusedSum(Posit32[],Quire).0._State\ := \Posit32::FusedSum(Posit32[],Quire).0._State_8\;
                            end if;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Quire Posit32::op_Explicit(Posit32).0._StateMachine\: process (\Clock\) 
        Variable \Quire Posit32::op_Explicit(Posit32).0._State\: \Quire Posit32::op_Explicit(Posit32).0._States\ := \Quire Posit32::op_Explicit(Posit32).0._State_0\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.x\: \Lombiq.Arithmetics.Posit32\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.this_2cf6f4dc9cc2c5c30dc9a398865472e185402e2a019e7ac16cc5146e4f812825\: \Lombiq.Arithmetics.Posit32\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_2cf6f4dc9cc2c5c30dc9a398865472e185402e2a019e7ac16cc5146e4f812825\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.0\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.objectced560230eaa29c09194274d79f0f04aeb95c7628d7ce6b644348e51440adb36\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.return.0\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.array\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
        Variable \Quire Posit32::op_Explicit(Posit32).0.this_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: \Lombiq.Arithmetics.Posit32\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.num_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.this_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: \Lombiq.Arithmetics.Posit32\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.bits_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.conditional963d17004b6788ad55358cce58986fa179ec1b5dc039dfede93d706448099e92_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.this_092f045227f64eda72b3fc95be3c3637705914add72214a343e55185cfa65c10_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: \Lombiq.Arithmetics.Posit32\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_092f045227f64eda72b3fc95be3c3637705914add72214a343e55185cfa65c10_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.1\: signed(63 downto 0) := to_signed(0, 64);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.2\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.bits_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.0\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.num_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.startingPosition_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.b_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.4\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.5\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.num_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.6\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.7\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.8\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.num2_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.9\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.10\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.11\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.12\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.13\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.14\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.15\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.16\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.17\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.18\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.conditionalf2eba7c459dd057c9270f346c2a9013399b4309fc21683746ef1be47061f03f1_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.19\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.num2_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.conditionalec88d618fdb8d955a353066f43af5ab5cc70c1913e02ecac14c3590c5ee9802e_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.this_21b5a692eb0046a4533a6168005ecc761e6f077932e1ccbe536f04342ca83a96_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: \Lombiq.Arithmetics.Posit32\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_21b5a692eb0046a4533a6168005ecc761e6f077932e1ccbe536f04342ca83a96_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.20\: signed(63 downto 0) := to_signed(0, 64);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.21\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.bits_0f83a95a96264a09c6a0ba9cb9c99ad3bd58dcf2757ca4c9081ded388086ca02_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_0f83a95a96264a09c6a0ba9cb9c99ad3bd58dcf2757ca4c9081ded388086ca02_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.1\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.22\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.bits_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.23\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.24\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.25\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.26\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.conditional7e2c70f465bbd6af6328e84460df8cc63262cd5e429e5f14f0c6d6c3620c3cea_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.27\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.this_fb93a852800b1e46e7592da171e65de7ddd0018d517ad2135ba24c2440a2f0e3_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: \Lombiq.Arithmetics.Posit32\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.bits_fb93a852800b1e46e7592da171e65de7ddd0018d517ad2135ba24c2440a2f0e3_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.index_fb93a852800b1e46e7592da171e65de7ddd0018d517ad2135ba24c2440a2f0e3_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_fb93a852800b1e46e7592da171e65de7ddd0018d517ad2135ba24c2440a2f0e3_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.28\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.29\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.quire\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.this_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\: \Lombiq.Arithmetics.Posit32\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.bits_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.conditional963d17004b6788ad55358cce58986fa179ec1b5dc039dfede93d706448099e92_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.this_092f045227f64eda72b3fc95be3c3637705914add72214a343e55185cfa65c10_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\: \Lombiq.Arithmetics.Posit32\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_092f045227f64eda72b3fc95be3c3637705914add72214a343e55185cfa65c10_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.30\: signed(63 downto 0) := to_signed(0, 64);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.31\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.bits_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.32\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.num_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.startingPosition_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.b_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.33\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.34\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.num_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.35\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.36\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.37\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.num2_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.38\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.39\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.40\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.41\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.42\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.43\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.44\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.45\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.46\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.47\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.conditionalf2eba7c459dd057c9270f346c2a9013399b4309fc21683746ef1be47061f03f1_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.48\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.this_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: \Lombiq.Arithmetics.Posit32\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: signed(15 downto 0) := to_signed(0, 16);
        Variable \Quire Posit32::op_Explicit(Posit32).0.regimeKValue_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: signed(7 downto 0) := to_signed(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.this_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: \Lombiq.Arithmetics.Posit32\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: signed(7 downto 0) := to_signed(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.num_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.conditional054ffdc2634715c514e630840f155e53d1c8ffe0be53ec06d4c21ba08ad2b716_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.this_7c713771ddbe04c4c2ff20ebfa1dae4044757c440fe5b46ea759182bcfb4b09b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: \Lombiq.Arithmetics.Posit32\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_7c713771ddbe04c4c2ff20ebfa1dae4044757c440fe5b46ea759182bcfb4b09b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.49\: signed(63 downto 0) := to_signed(0, 64);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.50\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.bits_6618db8f62e3464b32c8cc3e2209d7d35e6f677ff842c32f9130d90de0560ee2_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_6618db8f62e3464b32c8cc3e2209d7d35e6f677ff842c32f9130d90de0560ee2_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.3\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.51\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.bits_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.startingPosition_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.b_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.52\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.53\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.num_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.54\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.55\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.56\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.num2_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.57\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.58\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.59\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.60\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.61\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.62\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.63\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.conditional882cd98d817375e03765080fbf2e91fcc69740961af08057feb5bee6e57e0737_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: signed(7 downto 0) := to_signed(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.64\: signed(63 downto 0) := to_signed(0, 64);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.65\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.4\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.66\: signed(7 downto 0) := to_signed(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.conditional1aa95b35288eb627929161a1ee637479589960934567100c958634e64afb13de_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.67\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.this_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: \Lombiq.Arithmetics.Posit32\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.num_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.conditional880d0f3a8d33b2428fb4e8a62e4174f93b0cc01cc9b8d6d16563b7d2d4e90992_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.this_4d92f321cba6244b5bb71509cbad78bd467f0d9f83f5164197b9be70bc739dc2\: \Lombiq.Arithmetics.Posit32\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_4d92f321cba6244b5bb71509cbad78bd467f0d9f83f5164197b9be70bc739dc2\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.68\: signed(63 downto 0) := to_signed(0, 64);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.69\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.bits_c6f8839606b9f7c5e666e7f8d7c6eeb396a41e4838bd7ee0d04170e34ce7b814\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_c6f8839606b9f7c5e666e7f8d7c6eeb396a41e4838bd7ee0d04170e34ce7b814\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.5\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.70\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.b_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.this_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\: \Lombiq.Arithmetics.Posit32\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.bits_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.conditional85ca8d8893aa24483d9e74ed87417b722b6d33d6069def85ee5195c77759eab3_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.this_8ccfdac761d94cefabb354727c4eec638b4b892c15d704db2d4988c8e2e41cd8_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\: \Lombiq.Arithmetics.Posit32\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_8ccfdac761d94cefabb354727c4eec638b4b892c15d704db2d4988c8e2e41cd8_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.71\: signed(63 downto 0) := to_signed(0, 64);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.72\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.bits_3465d1fb5b2deaf339333582b5a596bf893ed003380b440bf76067c5451863a3_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_3465d1fb5b2deaf339333582b5a596bf893ed003380b440bf76067c5451863a3_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.6\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.73\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.bits_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.startingPosition_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.b_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.74\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.75\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.num_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.76\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.77\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.78\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.num2_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.79\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.80\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.81\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.82\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.83\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.84\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.85\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.86\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.87\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.conditional68bcd4673000ed90d5e5bddf9742548ff8843dd36c272b449a1de261af0ae5a9_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.88\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.89\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.90\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.91\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.92\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.93\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.94\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.this_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\: \Lombiq.Arithmetics.Posit32\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.bits_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.conditional963d17004b6788ad55358cce58986fa179ec1b5dc039dfede93d706448099e92_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.this_092f045227f64eda72b3fc95be3c3637705914add72214a343e55185cfa65c10_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\: \Lombiq.Arithmetics.Posit32\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_092f045227f64eda72b3fc95be3c3637705914add72214a343e55185cfa65c10_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.95\: signed(63 downto 0) := to_signed(0, 64);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.96\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.bits_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.7\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.97\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.num_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.startingPosition_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.b_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.98\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.99\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.num_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.100\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.101\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.102\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.num2_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.103\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.104\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.105\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.106\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.107\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.108\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.109\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.110\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.111\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.112\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.conditionalf2eba7c459dd057c9270f346c2a9013399b4309fc21683746ef1be47061f03f1_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.113\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.114\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.115\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.116\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.117\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.conditionala233560fe7dfff22c231bec46671f442fee11494dc774056e64d669ec36cdb00_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.118\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.119\: signed(63 downto 0) := to_signed(0, 64);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.120\: signed(15 downto 0) := to_signed(0, 16);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.121\: signed(63 downto 0) := to_signed(0, 64);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.122\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Posit32::op_Explicit(Posit32).0.return.1\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.this_5204dd194817ce0e22c54ac6e6fe7dc0a0e40352e5a5fed887c54294684dded0\: \Lombiq.Arithmetics.Posit32\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.return_5204dd194817ce0e22c54ac6e6fe7dc0a0e40352e5a5fed887c54294684dded0\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.123\: signed(63 downto 0) := to_signed(0, 64);
        Variable \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.124\: boolean := false;
        Variable \Quire Posit32::op_Explicit(Posit32).0.return.2\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire Posit32::op_Explicit(Posit32).0.return.3\: \Lombiq.Arithmetics.Quire\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Quire Posit32::op_Explicit(Posit32).0._Finished\ <= false;
                \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16).firstSegment.parameter.Out.0\ <= to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16)._Started.0\ <= false;
                \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\ <= to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ <= false;
                \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 64));
                \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= false;
                \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_OnesComplement(Quire)._Started.0\ <= false;
                \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32).right.parameter.Out.0\ <= to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32)._Started.0\ <= false;
                \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_0\;
                \Quire Posit32::op_Explicit(Posit32).0.return_2cf6f4dc9cc2c5c30dc9a398865472e185402e2a019e7ac16cc5146e4f812825\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.0\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.array\ := (others => to_unsigned(0, 64));
                \Quire Posit32::op_Explicit(Posit32).0.return_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.num_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.return_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.bits_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.conditional963d17004b6788ad55358cce58986fa179ec1b5dc039dfede93d706448099e92_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.return_092f045227f64eda72b3fc95be3c3637705914add72214a343e55185cfa65c10_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.1\ := to_signed(0, 64);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.2\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.bits_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.return_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.0\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.3\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.num_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.startingPosition_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.return_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.b_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.4\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.5\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.num_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.6\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.7\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.8\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.num2_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.9\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.10\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.11\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.12\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.13\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.14\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.15\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.16\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.17\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.18\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.conditionalf2eba7c459dd057c9270f346c2a9013399b4309fc21683746ef1be47061f03f1_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.19\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.num2_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.conditionalec88d618fdb8d955a353066f43af5ab5cc70c1913e02ecac14c3590c5ee9802e_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.return_21b5a692eb0046a4533a6168005ecc761e6f077932e1ccbe536f04342ca83a96_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.20\ := to_signed(0, 64);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.21\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.bits_0f83a95a96264a09c6a0ba9cb9c99ad3bd58dcf2757ca4c9081ded388086ca02_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.return_0f83a95a96264a09c6a0ba9cb9c99ad3bd58dcf2757ca4c9081ded388086ca02_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.1\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.22\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.bits_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.23\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.24\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.25\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.26\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.conditional7e2c70f465bbd6af6328e84460df8cc63262cd5e429e5f14f0c6d6c3620c3cea_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.27\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.bits_fb93a852800b1e46e7592da171e65de7ddd0018d517ad2135ba24c2440a2f0e3_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.index_fb93a852800b1e46e7592da171e65de7ddd0018d517ad2135ba24c2440a2f0e3_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(0, 16);
                \Quire Posit32::op_Explicit(Posit32).0.return_fb93a852800b1e46e7592da171e65de7ddd0018d517ad2135ba24c2440a2f0e3_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.28\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.29\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.return_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.bits_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.conditional963d17004b6788ad55358cce58986fa179ec1b5dc039dfede93d706448099e92_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.return_092f045227f64eda72b3fc95be3c3637705914add72214a343e55185cfa65c10_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.30\ := to_signed(0, 64);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.31\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.bits_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.return_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.2\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.32\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.num_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.startingPosition_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.return_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.b_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.33\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.34\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.num_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.35\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.36\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.37\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.num2_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.38\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.39\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.40\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.41\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.42\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.43\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.44\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.45\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.46\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.47\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.conditionalf2eba7c459dd057c9270f346c2a9013399b4309fc21683746ef1be47061f03f1_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.48\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.return_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_signed(0, 16);
                \Quire Posit32::op_Explicit(Posit32).0.regimeKValue_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_signed(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.return_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_signed(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.num_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.conditional054ffdc2634715c514e630840f155e53d1c8ffe0be53ec06d4c21ba08ad2b716_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.return_7c713771ddbe04c4c2ff20ebfa1dae4044757c440fe5b46ea759182bcfb4b09b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.49\ := to_signed(0, 64);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.50\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.bits_6618db8f62e3464b32c8cc3e2209d7d35e6f677ff842c32f9130d90de0560ee2_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.return_6618db8f62e3464b32c8cc3e2209d7d35e6f677ff842c32f9130d90de0560ee2_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.3\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.51\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.bits_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.startingPosition_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.return_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.b_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.52\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.53\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.num_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.54\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.55\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.56\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.num2_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.57\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.58\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.59\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.60\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.61\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.62\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.63\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.conditional882cd98d817375e03765080fbf2e91fcc69740961af08057feb5bee6e57e0737_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_signed(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.64\ := to_signed(0, 64);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.65\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.4\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.66\ := to_signed(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.conditional1aa95b35288eb627929161a1ee637479589960934567100c958634e64afb13de_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.67\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.return_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.num_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.conditional880d0f3a8d33b2428fb4e8a62e4174f93b0cc01cc9b8d6d16563b7d2d4e90992_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.return_4d92f321cba6244b5bb71509cbad78bd467f0d9f83f5164197b9be70bc739dc2\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.68\ := to_signed(0, 64);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.69\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.bits_c6f8839606b9f7c5e666e7f8d7c6eeb396a41e4838bd7ee0d04170e34ce7b814\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.return_c6f8839606b9f7c5e666e7f8d7c6eeb396a41e4838bd7ee0d04170e34ce7b814\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.5\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.70\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.b_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.return_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.bits_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.conditional85ca8d8893aa24483d9e74ed87417b722b6d33d6069def85ee5195c77759eab3_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.return_8ccfdac761d94cefabb354727c4eec638b4b892c15d704db2d4988c8e2e41cd8_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.71\ := to_signed(0, 64);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.72\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.bits_3465d1fb5b2deaf339333582b5a596bf893ed003380b440bf76067c5451863a3_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.return_3465d1fb5b2deaf339333582b5a596bf893ed003380b440bf76067c5451863a3_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.6\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.73\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.bits_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.startingPosition_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.return_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.b_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.74\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.75\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.num_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.76\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.77\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.78\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.num2_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.79\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.80\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.81\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.82\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.83\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.84\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.85\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.86\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.87\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.conditional68bcd4673000ed90d5e5bddf9742548ff8843dd36c272b449a1de261af0ae5a9_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.88\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.89\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.90\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.91\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.92\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.93\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.94\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.return_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.bits_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.conditional963d17004b6788ad55358cce58986fa179ec1b5dc039dfede93d706448099e92_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.return_092f045227f64eda72b3fc95be3c3637705914add72214a343e55185cfa65c10_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.95\ := to_signed(0, 64);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.96\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.bits_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.return_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.7\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.97\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.num_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.startingPosition_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.return_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.b_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.98\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.99\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.num_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.100\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.101\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.102\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.num2_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.103\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.104\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.105\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.106\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.107\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.108\ := to_unsigned(0, 8);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.109\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.110\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.111\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.112\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.conditionalf2eba7c459dd057c9270f346c2a9013399b4309fc21683746ef1be47061f03f1_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.113\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.114\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.115\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.116\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.117\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.conditionala233560fe7dfff22c231bec46671f442fee11494dc774056e64d669ec36cdb00_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_unsigned(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.118\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.119\ := to_signed(0, 64);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.120\ := to_signed(0, 16);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.121\ := to_signed(0, 64);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.122\ := to_signed(0, 32);
                \Quire Posit32::op_Explicit(Posit32).0.return_5204dd194817ce0e22c54ac6e6fe7dc0a0e40352e5a5fed887c54294684dded0\ := false;
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.123\ := to_signed(0, 64);
                \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.124\ := false;
            else 
                case \Quire Posit32::op_Explicit(Posit32).0._State\ is 
                    when \Quire Posit32::op_Explicit(Posit32).0._State_0\ => 
                        
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._Started\ = true) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_2\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_1\ => 
                        
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._Started\ = true) then 
                            \Quire Posit32::op_Explicit(Posit32).0._Finished\ <= true;
                        else 
                            \Quire Posit32::op_Explicit(Posit32).0._Finished\ <= false;
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_0\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_2\ => 
                        \Quire Posit32::op_Explicit(Posit32).0.x\ := \Quire Posit32::op_Explicit(Posit32).0.x.parameter.In\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.this_2cf6f4dc9cc2c5c30dc9a398865472e185402e2a019e7ac16cc5146e4f812825\ := \Quire Posit32::op_Explicit(Posit32).0.x\;
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.0\ := \Quire Posit32::op_Explicit(Posit32).0.this_2cf6f4dc9cc2c5c30dc9a398865472e185402e2a019e7ac16cc5146e4f812825\.\PositBits\ = "10000000000000000000000000000000";
                        \Quire Posit32::op_Explicit(Posit32).0.return_2cf6f4dc9cc2c5c30dc9a398865472e185402e2a019e7ac16cc5146e4f812825\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.0\;
                        
                        
                        
                        
                        
                        
                        

                        
                        
                        

                        if (\Quire Posit32::op_Explicit(Posit32).0.return_2cf6f4dc9cc2c5c30dc9a398865472e185402e2a019e7ac16cc5146e4f812825\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_5\;
                        else 
                            
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_4\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_3\ => 
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.b_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.return_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\;
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.this_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := \Quire Posit32::op_Explicit(Posit32).0.this_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.this_092f045227f64eda72b3fc95be3c3637705914add72214a343e55185cfa65c10_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := \Quire Posit32::op_Explicit(Posit32).0.this_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\;
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.95\ := signed(SmartResize(\Quire Posit32::op_Explicit(Posit32).0.this_092f045227f64eda72b3fc95be3c3637705914add72214a343e55185cfa65c10_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\.\PositBits\ and "10000000000000000000000000000000", 64));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.96\ := signed(SmartResize(((\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.95\)), 64)) = to_signed(0, 64);
                        \Quire Posit32::op_Explicit(Posit32).0.return_092f045227f64eda72b3fc95be3c3637705914add72214a343e55185cfa65c10_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.96\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        

                        
                        
                        
                        

                        if (\Quire Posit32::op_Explicit(Posit32).0.return_092f045227f64eda72b3fc95be3c3637705914add72214a343e55185cfa65c10_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_74\;
                        else 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_75\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_4\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.array\ := (others => to_unsigned(0, 64));
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.this_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.x\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.this_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.this_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.this_092f045227f64eda72b3fc95be3c3637705914add72214a343e55185cfa65c10_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.this_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\;
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.1\ := signed(SmartResize(\Quire Posit32::op_Explicit(Posit32).0.this_092f045227f64eda72b3fc95be3c3637705914add72214a343e55185cfa65c10_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\.\PositBits\ and "10000000000000000000000000000000", 64));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.2\ := signed(SmartResize(((\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.1\)), 64)) = to_signed(0, 64);
                        \Quire Posit32::op_Explicit(Posit32).0.return_092f045227f64eda72b3fc95be3c3637705914add72214a343e55185cfa65c10_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.2\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        

                        
                        
                        
                        

                        if (\Quire Posit32::op_Explicit(Posit32).0.return_092f045227f64eda72b3fc95be3c3637705914add72214a343e55185cfa65c10_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_9\;
                        else 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_10\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_5\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.objectced560230eaa29c09194274d79f0f04aeb95c7628d7ce6b644348e51440adb36\.\IsNull\ := false;
                        \Quire Posit32::op_Explicit(Posit32).0.objectced560230eaa29c09194274d79f0f04aeb95c7628d7ce6b644348e51440adb36\.\Size\ := to_unsigned(0, 16);
                        \Quire Posit32::op_Explicit(Posit32).0.objectced560230eaa29c09194274d79f0f04aeb95c7628d7ce6b644348e51440adb36\.\SegmentCount\ := to_unsigned(0, 16);
                        \Quire Posit32::op_Explicit(Posit32).0.objectced560230eaa29c09194274d79f0f04aeb95c7628d7ce6b644348e51440adb36\.\Segments\ := (others => to_unsigned(0, 64));
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16).this.parameter.Out.0\ <= \Quire Posit32::op_Explicit(Posit32).0.objectced560230eaa29c09194274d79f0f04aeb95c7628d7ce6b644348e51440adb36\;
                        \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16).firstSegment.parameter.Out.0\ <= to_unsigned(1, 32);
                        \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16).size.parameter.Out.0\ <= SmartResize(unsigned(to_signed(512, 32)), 16);
                        \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16)._Started.0\ <= true;
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_6\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_6\ => 
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16)._Started.0\ = \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16)._Finished.0\) then 
                            \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16)._Started.0\ <= false;
                            \Quire Posit32::op_Explicit(Posit32).0.objectced560230eaa29c09194274d79f0f04aeb95c7628d7ce6b644348e51440adb36\ := \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16).this.parameter.In.0\;
                            
                            
                            
                            
                            \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.Out.0\ <= \Quire Posit32::op_Explicit(Posit32).0.objectced560230eaa29c09194274d79f0f04aeb95c7628d7ce6b644348e51440adb36\;
                            \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\ <= to_signed(511, 32);
                            \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ <= true;
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_7\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_7\ => 
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ = \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\) then 
                            \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ <= false;
                            \Quire Posit32::op_Explicit(Posit32).0.return.0\ := \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).return.0\;
                            \Quire Posit32::op_Explicit(Posit32).0.objectced560230eaa29c09194274d79f0f04aeb95c7628d7ce6b644348e51440adb36\ := \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.In.0\;
                            \Quire Posit32::op_Explicit(Posit32).0.return\ <= \Quire Posit32::op_Explicit(Posit32).0.return.0\;
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_1\;
                            
                            if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_7\) then 
                                \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_4\;
                            end if;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_8\ => 
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.bits_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := (\Quire Posit32::op_Explicit(Posit32).0.conditional963d17004b6788ad55358cce58986fa179ec1b5dc039dfede93d706448099e92_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.bits_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\;
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.startingPosition_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := SmartResize(unsigned(to_signed(31, 32)), 8);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.b_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := SmartResize(unsigned(to_signed(1, 32)), 8);
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.4\ := to_signed(32, 32) - signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.startingPosition_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\), 32));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.5\ := shift_left(\Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\, to_integer(unsigned(SmartResize(\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.4\, 5))));
                        \Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.5\;
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_11\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_9\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditional963d17004b6788ad55358cce58986fa179ec1b5dc039dfede93d706448099e92_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.this_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\.\PositBits\;
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_9\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_8\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_10\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.bits_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.this_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\.\PositBits\;
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.0\ := not(\Quire Posit32::op_Explicit(Posit32).0.bits_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\);
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.3\ := SmartResize(unsigned(signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.0\), 64)) + to_signed(1, 64)), 32);
                        \Quire Posit32::op_Explicit(Posit32).0.return_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.3\);
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditional963d17004b6788ad55358cce58986fa179ec1b5dc039dfede93d706448099e92_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.return_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\;
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_10\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_8\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_11\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.6\ := shift_right(\Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\, to_integer(unsigned(SmartResize(to_signed(31, 32), 5) and "11111")));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.7\ := (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.6\) and to_unsigned(1, 32);
                        \Quire Posit32::op_Explicit(Posit32).0.num_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.7\;
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.8\ := shift_left(\Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\, to_integer(unsigned(SmartResize(to_signed(1, 32), 5))));
                        \Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.8\;
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.num2_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_signed(0, 32);
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_12\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_12\ => 
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.9\ := (\Quire Posit32::op_Explicit(Posit32).0.num2_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\) < signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.startingPosition_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\), 32));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.10\ := shift_right(\Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\, to_integer(unsigned(SmartResize(to_signed(31, 32), 5) and "11111")));
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_14\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_13\ => 
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.return_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.b_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\;
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.16\ := signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.return_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\), 32)) + to_signed(2, 32);
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.17\ := SmartResize(\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.16\ + to_signed(2, 32), 32);
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_16\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_14\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.11\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.10\ = \Quire Posit32::op_Explicit(Posit32).0.num_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\;
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.12\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.9\ and \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.11\;
                        if (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.12\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.13\ := shift_left(\Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\, to_integer(unsigned(SmartResize(to_signed(1, 32), 5))));
                            \Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.13\;
                            
                            
                            
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_15\;
                        else 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_13\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_15\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.14\ := SmartResize(unsigned(signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.b_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\), 32)) + to_signed(1, 32)), 8);
                        \Quire Posit32::op_Explicit(Posit32).0.b_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.14\);
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.15\ := \Quire Posit32::op_Explicit(Posit32).0.num2_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ + to_signed(1, 32);
                        \Quire Posit32::op_Explicit(Posit32).0.num2_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.15\;
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_15\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_12\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_16\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.18\ := to_signed(32, 32) - (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.17\);
                        \Quire Posit32::op_Explicit(Posit32).0.num_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.18\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.19\ := \Quire Posit32::op_Explicit(Posit32).0.num_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ > to_signed(0, 32);

                        
                        
                        
                        

                        if ((\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.19\)) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_18\;
                        else 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_19\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_17\ => 
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.return_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.conditionalf2eba7c459dd057c9270f346c2a9013399b4309fc21683746ef1be47061f03f1_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\;
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.num_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.return_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.this_21b5a692eb0046a4533a6168005ecc761e6f077932e1ccbe536f04342ca83a96_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.this_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\;
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.20\ := signed(SmartResize(\Quire Posit32::op_Explicit(Posit32).0.this_21b5a692eb0046a4533a6168005ecc761e6f077932e1ccbe536f04342ca83a96_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\.\PositBits\ and "10000000000000000000000000000000", 64));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.21\ := signed(SmartResize(((\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.20\)), 64)) = to_signed(0, 64);
                        \Quire Posit32::op_Explicit(Posit32).0.return_21b5a692eb0046a4533a6168005ecc761e6f077932e1ccbe536f04342ca83a96_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.21\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        

                        
                        
                        
                        

                        if (\Quire Posit32::op_Explicit(Posit32).0.return_21b5a692eb0046a4533a6168005ecc761e6f077932e1ccbe536f04342ca83a96_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_21\;
                        else 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_22\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_18\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditionalf2eba7c459dd057c9270f346c2a9013399b4309fc21683746ef1be47061f03f1_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := (unsigned(\Quire Posit32::op_Explicit(Posit32).0.num_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\));
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_18\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_17\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_19\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditionalf2eba7c459dd057c9270f346c2a9013399b4309fc21683746ef1be47061f03f1_c19fcd84e7300e48def129d35eb60d7e89695194c445b7224655f2d93aee9a18_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(0, 32);
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_19\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_17\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_20\ => 
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.num2_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := (\Quire Posit32::op_Explicit(Posit32).0.conditionalec88d618fdb8d955a353066f43af5ab5cc70c1913e02ecac14c3590c5ee9802e_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\);
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.23\ := SmartResize(to_signed(32, 64) - signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.num_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\), 64)), 32);
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.24\ := shift_left(\Quire Posit32::op_Explicit(Posit32).0.num2_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\, to_integer(unsigned(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.23\), 5))));
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_23\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_21\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditionalec88d618fdb8d955a353066f43af5ab5cc70c1913e02ecac14c3590c5ee9802e_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.this_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\.\PositBits\;
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_21\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_20\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_22\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.bits_0f83a95a96264a09c6a0ba9cb9c99ad3bd58dcf2757ca4c9081ded388086ca02_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.this_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\.\PositBits\;
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.1\ := not(\Quire Posit32::op_Explicit(Posit32).0.bits_0f83a95a96264a09c6a0ba9cb9c99ad3bd58dcf2757ca4c9081ded388086ca02_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\);
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.22\ := SmartResize(unsigned(signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.1\), 64)) + to_signed(1, 64)), 32);
                        \Quire Posit32::op_Explicit(Posit32).0.return_0f83a95a96264a09c6a0ba9cb9c99ad3bd58dcf2757ca4c9081ded388086ca02_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.22\);
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditionalec88d618fdb8d955a353066f43af5ab5cc70c1913e02ecac14c3590c5ee9802e_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.return_0f83a95a96264a09c6a0ba9cb9c99ad3bd58dcf2757ca4c9081ded388086ca02_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\;
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_22\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_20\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_23\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.25\ := SmartResize(to_signed(32, 64) - signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.num_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\), 64)), 32);
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_24\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_24\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.26\ := shift_right(\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.24\, to_integer(unsigned(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.25\), 5) and "11111")));
                        \Quire Posit32::op_Explicit(Posit32).0.bits_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.26\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_25\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_25\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.27\ := signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.num_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\), 64)) = to_signed(0, 64);

                        
                        
                        
                        

                        if ((\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.27\)) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_27\;
                        else 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_28\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_26\ => 
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.return_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.conditional7e2c70f465bbd6af6328e84460df8cc63262cd5e429e5f14f0c6d6c3620c3cea_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\;
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.array\(to_integer(to_signed(0, 32))) := SmartResize(\Quire Posit32::op_Explicit(Posit32).0.return_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\, 64);
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.quire\.\IsNull\ := false;
                        \Quire Posit32::op_Explicit(Posit32).0.quire\.\Size\ := to_unsigned(0, 16);
                        \Quire Posit32::op_Explicit(Posit32).0.quire\.\SegmentCount\ := to_unsigned(0, 16);
                        \Quire Posit32::op_Explicit(Posit32).0.quire\.\Segments\ := (others => to_unsigned(0, 64));
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\ <= \Quire Posit32::op_Explicit(Posit32).0.quire\;
                        \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\ <= \Quire Posit32::op_Explicit(Posit32).0.array\;
                        \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\ <= SmartResize(unsigned(to_signed(0, 32)), 16);
                        \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= true;
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_29\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_27\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditional7e2c70f465bbd6af6328e84460df8cc63262cd5e429e5f14f0c6d6c3620c3cea_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := to_unsigned(1, 32);
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_27\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_26\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_28\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.this_fb93a852800b1e46e7592da171e65de7ddd0018d517ad2135ba24c2440a2f0e3_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.this_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\;
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.bits_fb93a852800b1e46e7592da171e65de7ddd0018d517ad2135ba24c2440a2f0e3_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.bits_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\;
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.index_fb93a852800b1e46e7592da171e65de7ddd0018d517ad2135ba24c2440a2f0e3_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := SmartResize(\Quire Posit32::op_Explicit(Posit32).0.num_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\, 16);
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.28\ := unsigned(shift_left(to_signed(1, 32), to_integer(unsigned(SmartResize(signed(SmartResize(\Quire Posit32::op_Explicit(Posit32).0.index_fb93a852800b1e46e7592da171e65de7ddd0018d517ad2135ba24c2440a2f0e3_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\, 32)), 5)))));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.29\ := \Quire Posit32::op_Explicit(Posit32).0.bits_fb93a852800b1e46e7592da171e65de7ddd0018d517ad2135ba24c2440a2f0e3_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ or (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.28\);
                        \Quire Posit32::op_Explicit(Posit32).0.return_fb93a852800b1e46e7592da171e65de7ddd0018d517ad2135ba24c2440a2f0e3_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.29\;
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditional7e2c70f465bbd6af6328e84460df8cc63262cd5e429e5f14f0c6d6c3620c3cea_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\ := \Quire Posit32::op_Explicit(Posit32).0.return_fb93a852800b1e46e7592da171e65de7ddd0018d517ad2135ba24c2440a2f0e3_310be957880a463aabf2b9e3fe034bc10c979fe352d91dac9b2227df64d3429d\;
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_28\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_26\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_29\ => 
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ = \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\) then 
                            \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= false;
                            \Quire Posit32::op_Explicit(Posit32).0.quire\ := \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\;
                            \Quire Posit32::op_Explicit(Posit32).0.array\ := \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\;
                            
                            
                            
                            
                            
                            
                            \Quire Posit32::op_Explicit(Posit32).0.this_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := \Quire Posit32::op_Explicit(Posit32).0.x\;
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Posit32::op_Explicit(Posit32).0.this_092f045227f64eda72b3fc95be3c3637705914add72214a343e55185cfa65c10_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := \Quire Posit32::op_Explicit(Posit32).0.this_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\;
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.30\ := signed(SmartResize(\Quire Posit32::op_Explicit(Posit32).0.this_092f045227f64eda72b3fc95be3c3637705914add72214a343e55185cfa65c10_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\.\PositBits\ and "10000000000000000000000000000000", 64));
                            \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.31\ := signed(SmartResize(((\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.30\)), 64)) = to_signed(0, 64);
                            \Quire Posit32::op_Explicit(Posit32).0.return_092f045227f64eda72b3fc95be3c3637705914add72214a343e55185cfa65c10_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.31\;
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            

                            
                            
                            
                            

                            if (\Quire Posit32::op_Explicit(Posit32).0.return_092f045227f64eda72b3fc95be3c3637705914add72214a343e55185cfa65c10_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\) then 
                                \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_31\;
                            else 
                                \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_32\;
                            end if;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_30\ => 
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.bits_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := (\Quire Posit32::op_Explicit(Posit32).0.conditional963d17004b6788ad55358cce58986fa179ec1b5dc039dfede93d706448099e92_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := \Quire Posit32::op_Explicit(Posit32).0.bits_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\;
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.startingPosition_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := SmartResize(unsigned(to_signed(31, 32)), 8);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.b_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := SmartResize(unsigned(to_signed(1, 32)), 8);
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.33\ := to_signed(32, 32) - signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.startingPosition_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\), 32));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.34\ := shift_left(\Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\, to_integer(unsigned(SmartResize(\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.33\, 5))));
                        \Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.34\;
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_33\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_31\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditional963d17004b6788ad55358cce58986fa179ec1b5dc039dfede93d706448099e92_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := \Quire Posit32::op_Explicit(Posit32).0.this_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\.\PositBits\;
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_31\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_30\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_32\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.bits_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := \Quire Posit32::op_Explicit(Posit32).0.this_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\.\PositBits\;
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.2\ := not(\Quire Posit32::op_Explicit(Posit32).0.bits_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\);
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.32\ := SmartResize(unsigned(signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.2\), 64)) + to_signed(1, 64)), 32);
                        \Quire Posit32::op_Explicit(Posit32).0.return_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.32\);
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditional963d17004b6788ad55358cce58986fa179ec1b5dc039dfede93d706448099e92_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := \Quire Posit32::op_Explicit(Posit32).0.return_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\;
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_32\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_30\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_33\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.35\ := shift_right(\Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\, to_integer(unsigned(SmartResize(to_signed(31, 32), 5) and "11111")));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.36\ := (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.35\) and to_unsigned(1, 32);
                        \Quire Posit32::op_Explicit(Posit32).0.num_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.36\;
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.37\ := shift_left(\Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\, to_integer(unsigned(SmartResize(to_signed(1, 32), 5))));
                        \Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.37\;
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.num2_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := to_signed(0, 32);
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_34\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_34\ => 
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.38\ := (\Quire Posit32::op_Explicit(Posit32).0.num2_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\) < signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.startingPosition_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\), 32));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.39\ := shift_right(\Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\, to_integer(unsigned(SmartResize(to_signed(31, 32), 5) and "11111")));
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_36\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_35\ => 
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.return_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := \Quire Posit32::op_Explicit(Posit32).0.b_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\;
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.45\ := signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.return_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\), 32)) + to_signed(2, 32);
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.46\ := SmartResize(\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.45\ + to_signed(2, 32), 32);
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_38\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_36\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.40\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.39\ = \Quire Posit32::op_Explicit(Posit32).0.num_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\;
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.41\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.38\ and \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.40\;
                        if (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.41\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.42\ := shift_left(\Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\, to_integer(unsigned(SmartResize(to_signed(1, 32), 5))));
                            \Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.42\;
                            
                            
                            
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_37\;
                        else 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_35\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_37\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.43\ := SmartResize(unsigned(signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.b_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\), 32)) + to_signed(1, 32)), 8);
                        \Quire Posit32::op_Explicit(Posit32).0.b_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.43\);
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.44\ := \Quire Posit32::op_Explicit(Posit32).0.num2_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ + to_signed(1, 32);
                        \Quire Posit32::op_Explicit(Posit32).0.num2_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.44\;
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_37\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_34\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_38\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.47\ := to_signed(32, 32) - (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.46\);
                        \Quire Posit32::op_Explicit(Posit32).0.num_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.47\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.48\ := \Quire Posit32::op_Explicit(Posit32).0.num_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ > to_signed(0, 32);

                        
                        
                        
                        

                        if ((\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.48\)) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_40\;
                        else 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_41\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_39\ => 
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.return_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := \Quire Posit32::op_Explicit(Posit32).0.conditionalf2eba7c459dd057c9270f346c2a9013399b4309fc21683746ef1be47061f03f1_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\;
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.this_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.x\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.this_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.this_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.this_7c713771ddbe04c4c2ff20ebfa1dae4044757c440fe5b46ea759182bcfb4b09b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.this_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\;
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.49\ := signed(SmartResize(\Quire Posit32::op_Explicit(Posit32).0.this_7c713771ddbe04c4c2ff20ebfa1dae4044757c440fe5b46ea759182bcfb4b09b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\.\PositBits\ and "10000000000000000000000000000000", 64));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.50\ := signed(SmartResize(((\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.49\)), 64)) = to_signed(0, 64);
                        \Quire Posit32::op_Explicit(Posit32).0.return_7c713771ddbe04c4c2ff20ebfa1dae4044757c440fe5b46ea759182bcfb4b09b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.50\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        

                        
                        
                        
                        

                        if (\Quire Posit32::op_Explicit(Posit32).0.return_7c713771ddbe04c4c2ff20ebfa1dae4044757c440fe5b46ea759182bcfb4b09b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_43\;
                        else 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_44\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_40\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditionalf2eba7c459dd057c9270f346c2a9013399b4309fc21683746ef1be47061f03f1_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := (unsigned(\Quire Posit32::op_Explicit(Posit32).0.num_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\));
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_40\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_39\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_41\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditionalf2eba7c459dd057c9270f346c2a9013399b4309fc21683746ef1be47061f03f1_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\ := to_unsigned(0, 32);
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_41\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_39\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_42\ => 
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.num_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := (\Quire Posit32::op_Explicit(Posit32).0.conditional054ffdc2634715c514e630840f155e53d1c8ffe0be53ec06d4c21ba08ad2b716_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.bits_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.num_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\;
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.startingPosition_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := SmartResize(unsigned(to_signed(31, 32)), 8);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.b_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := SmartResize(unsigned(to_signed(1, 32)), 8);
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.52\ := to_signed(32, 32) - signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.startingPosition_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\), 32));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.53\ := shift_left(\Quire Posit32::op_Explicit(Posit32).0.bits_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\, to_integer(unsigned(SmartResize(\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.52\, 5))));
                        \Quire Posit32::op_Explicit(Posit32).0.bits_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.53\;
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_45\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_43\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditional054ffdc2634715c514e630840f155e53d1c8ffe0be53ec06d4c21ba08ad2b716_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.this_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\.\PositBits\;
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_43\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_42\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_44\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.bits_6618db8f62e3464b32c8cc3e2209d7d35e6f677ff842c32f9130d90de0560ee2_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.this_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\.\PositBits\;
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.3\ := not(\Quire Posit32::op_Explicit(Posit32).0.bits_6618db8f62e3464b32c8cc3e2209d7d35e6f677ff842c32f9130d90de0560ee2_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\);
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.51\ := SmartResize(unsigned(signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.3\), 64)) + to_signed(1, 64)), 32);
                        \Quire Posit32::op_Explicit(Posit32).0.return_6618db8f62e3464b32c8cc3e2209d7d35e6f677ff842c32f9130d90de0560ee2_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.51\);
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditional054ffdc2634715c514e630840f155e53d1c8ffe0be53ec06d4c21ba08ad2b716_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.return_6618db8f62e3464b32c8cc3e2209d7d35e6f677ff842c32f9130d90de0560ee2_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\;
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_44\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_42\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_45\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.54\ := shift_right(\Quire Posit32::op_Explicit(Posit32).0.bits_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\, to_integer(unsigned(SmartResize(to_signed(31, 32), 5) and "11111")));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.55\ := (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.54\) and to_unsigned(1, 32);
                        \Quire Posit32::op_Explicit(Posit32).0.num_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.55\;
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.56\ := shift_left(\Quire Posit32::op_Explicit(Posit32).0.bits_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\, to_integer(unsigned(SmartResize(to_signed(1, 32), 5))));
                        \Quire Posit32::op_Explicit(Posit32).0.bits_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.56\;
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.num2_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_signed(0, 32);
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_46\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_46\ => 
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.57\ := (\Quire Posit32::op_Explicit(Posit32).0.num2_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\) < signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.startingPosition_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\), 32));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.58\ := shift_right(\Quire Posit32::op_Explicit(Posit32).0.bits_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\, to_integer(unsigned(SmartResize(to_signed(31, 32), 5) and "11111")));
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_48\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_47\ => 
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.return_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.b_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\;
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.return_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.64\ := signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.num_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\), 64)) and to_signed(1073741824, 64);
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.65\ := (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.64\) = to_signed(0, 64);

                        
                        
                        
                        

                        if ((\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.65\)) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_51\;
                        else 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_52\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_48\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.59\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.58\ = \Quire Posit32::op_Explicit(Posit32).0.num_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\;
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.60\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.57\ and \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.59\;
                        if (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.60\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.61\ := shift_left(\Quire Posit32::op_Explicit(Posit32).0.bits_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\, to_integer(unsigned(SmartResize(to_signed(1, 32), 5))));
                            \Quire Posit32::op_Explicit(Posit32).0.bits_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.61\;
                            
                            
                            
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_49\;
                        else 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_47\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_49\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.62\ := SmartResize(unsigned(signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.b_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\), 32)) + to_signed(1, 32)), 8);
                        \Quire Posit32::op_Explicit(Posit32).0.b_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.62\);
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.63\ := \Quire Posit32::op_Explicit(Posit32).0.num2_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ + to_signed(1, 32);
                        \Quire Posit32::op_Explicit(Posit32).0.num2_99370110dae22db8631ca471eb437acc86c558e498739532bd9c0197bd7b376b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.63\;
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_49\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_46\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_50\ => 
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.return_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.conditional882cd98d817375e03765080fbf2e91fcc69740961af08057feb5bee6e57e0737_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\;
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.regimeKValue_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.return_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.67\ := SmartResize((\Quire Posit32::op_Explicit(Posit32).0.regimeKValue_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\), 32) /= to_signed(-31, 32);

                        
                        
                        
                        

                        if ((\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.67\)) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_54\;
                        else 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_90\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_51\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.4\ := -signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\), 32));
                        \Quire Posit32::op_Explicit(Posit32).0.conditional882cd98d817375e03765080fbf2e91fcc69740961af08057feb5bee6e57e0737_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := (SmartResize((\Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.4\), 8));
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_51\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_50\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_52\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.66\ := SmartResize(signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.b_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\), 32)) - to_signed(1, 32), 8);
                        \Quire Posit32::op_Explicit(Posit32).0.conditional882cd98d817375e03765080fbf2e91fcc69740961af08057feb5bee6e57e0737_832c1453bf6766412ab7d49a3bfbb4a30fb5f9d2e99fd33b1e1f82b95af141f7_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := ((\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.66\));
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_52\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_50\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_53\ => 
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.return_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := SmartResize((\Quire Posit32::op_Explicit(Posit32).0.conditional1aa95b35288eb627929161a1ee637479589960934567100c958634e64afb13de_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\), 16);
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.121\ := to_signed(240, 64) - signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.return_8dfbaed5965e93c29818d159b1ad2555bb8b028790c39ebb33911ab61c042d02\), 64));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.122\ := SmartResize(\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.121\ + SmartResize((\Quire Posit32::op_Explicit(Posit32).0.return_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\), 64), 32);
                        
                        \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.Out.0\ <= \Quire Posit32::op_Explicit(Posit32).0.quire\;
                        \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\ <= (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.122\);
                        \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ <= true;
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_91\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_54\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.this_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.this_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.this_4d92f321cba6244b5bb71509cbad78bd467f0d9f83f5164197b9be70bc739dc2\ := \Quire Posit32::op_Explicit(Posit32).0.this_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\;
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.68\ := signed(SmartResize(\Quire Posit32::op_Explicit(Posit32).0.this_4d92f321cba6244b5bb71509cbad78bd467f0d9f83f5164197b9be70bc739dc2\.\PositBits\ and "10000000000000000000000000000000", 64));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.69\ := signed(SmartResize(((\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.68\)), 64)) = to_signed(0, 64);
                        \Quire Posit32::op_Explicit(Posit32).0.return_4d92f321cba6244b5bb71509cbad78bd467f0d9f83f5164197b9be70bc739dc2\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.69\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        

                        
                        
                        
                        

                        if (\Quire Posit32::op_Explicit(Posit32).0.return_4d92f321cba6244b5bb71509cbad78bd467f0d9f83f5164197b9be70bc739dc2\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_56\;
                        else 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_57\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_55\ => 
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.num_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := (\Quire Posit32::op_Explicit(Posit32).0.conditional880d0f3a8d33b2428fb4e8a62e4174f93b0cc01cc9b8d6d16563b7d2d4e90992_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.this_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := \Quire Posit32::op_Explicit(Posit32).0.this_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.this_8ccfdac761d94cefabb354727c4eec638b4b892c15d704db2d4988c8e2e41cd8_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := \Quire Posit32::op_Explicit(Posit32).0.this_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\;
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.71\ := signed(SmartResize(\Quire Posit32::op_Explicit(Posit32).0.this_8ccfdac761d94cefabb354727c4eec638b4b892c15d704db2d4988c8e2e41cd8_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\.\PositBits\ and "10000000000000000000000000000000", 64));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.72\ := signed(SmartResize(((\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.71\)), 64)) = to_signed(0, 64);
                        \Quire Posit32::op_Explicit(Posit32).0.return_8ccfdac761d94cefabb354727c4eec638b4b892c15d704db2d4988c8e2e41cd8_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.72\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        

                        
                        
                        
                        

                        if (\Quire Posit32::op_Explicit(Posit32).0.return_8ccfdac761d94cefabb354727c4eec638b4b892c15d704db2d4988c8e2e41cd8_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_59\;
                        else 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_60\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_56\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditional880d0f3a8d33b2428fb4e8a62e4174f93b0cc01cc9b8d6d16563b7d2d4e90992_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.this_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\.\PositBits\;
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_56\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_55\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_57\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.bits_c6f8839606b9f7c5e666e7f8d7c6eeb396a41e4838bd7ee0d04170e34ce7b814\ := \Quire Posit32::op_Explicit(Posit32).0.this_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\.\PositBits\;
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.5\ := not(\Quire Posit32::op_Explicit(Posit32).0.bits_c6f8839606b9f7c5e666e7f8d7c6eeb396a41e4838bd7ee0d04170e34ce7b814\);
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.70\ := SmartResize(unsigned(signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.5\), 64)) + to_signed(1, 64)), 32);
                        \Quire Posit32::op_Explicit(Posit32).0.return_c6f8839606b9f7c5e666e7f8d7c6eeb396a41e4838bd7ee0d04170e34ce7b814\ := (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.70\);
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditional880d0f3a8d33b2428fb4e8a62e4174f93b0cc01cc9b8d6d16563b7d2d4e90992_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.return_c6f8839606b9f7c5e666e7f8d7c6eeb396a41e4838bd7ee0d04170e34ce7b814\;
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_57\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_55\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_58\ => 
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.bits_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := (\Quire Posit32::op_Explicit(Posit32).0.conditional85ca8d8893aa24483d9e74ed87417b722b6d33d6069def85ee5195c77759eab3_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.bits_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := \Quire Posit32::op_Explicit(Posit32).0.bits_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\;
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.startingPosition_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := SmartResize(unsigned(to_signed(31, 32)), 8);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.b_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := SmartResize(unsigned(to_signed(1, 32)), 8);
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.74\ := to_signed(32, 32) - signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.startingPosition_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\), 32));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.75\ := shift_left(\Quire Posit32::op_Explicit(Posit32).0.bits_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\, to_integer(unsigned(SmartResize(\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.74\, 5))));
                        \Quire Posit32::op_Explicit(Posit32).0.bits_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.75\;
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_61\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_59\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditional85ca8d8893aa24483d9e74ed87417b722b6d33d6069def85ee5195c77759eab3_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := \Quire Posit32::op_Explicit(Posit32).0.this_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\.\PositBits\;
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_59\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_58\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_60\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.bits_3465d1fb5b2deaf339333582b5a596bf893ed003380b440bf76067c5451863a3_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := \Quire Posit32::op_Explicit(Posit32).0.this_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\.\PositBits\;
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.6\ := not(\Quire Posit32::op_Explicit(Posit32).0.bits_3465d1fb5b2deaf339333582b5a596bf893ed003380b440bf76067c5451863a3_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\);
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.73\ := SmartResize(unsigned(signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.6\), 64)) + to_signed(1, 64)), 32);
                        \Quire Posit32::op_Explicit(Posit32).0.return_3465d1fb5b2deaf339333582b5a596bf893ed003380b440bf76067c5451863a3_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.73\);
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditional85ca8d8893aa24483d9e74ed87417b722b6d33d6069def85ee5195c77759eab3_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := \Quire Posit32::op_Explicit(Posit32).0.return_3465d1fb5b2deaf339333582b5a596bf893ed003380b440bf76067c5451863a3_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\;
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_60\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_58\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_61\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.76\ := shift_right(\Quire Posit32::op_Explicit(Posit32).0.bits_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\, to_integer(unsigned(SmartResize(to_signed(31, 32), 5) and "11111")));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.77\ := (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.76\) and to_unsigned(1, 32);
                        \Quire Posit32::op_Explicit(Posit32).0.num_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.77\;
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.78\ := shift_left(\Quire Posit32::op_Explicit(Posit32).0.bits_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\, to_integer(unsigned(SmartResize(to_signed(1, 32), 5))));
                        \Quire Posit32::op_Explicit(Posit32).0.bits_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.78\;
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.num2_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := to_signed(0, 32);
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_62\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_62\ => 
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.79\ := (\Quire Posit32::op_Explicit(Posit32).0.num2_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\) < signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.startingPosition_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\), 32));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.80\ := shift_right(\Quire Posit32::op_Explicit(Posit32).0.bits_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\, to_integer(unsigned(SmartResize(to_signed(31, 32), 5) and "11111")));
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_64\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_63\ => 
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.return_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := \Quire Posit32::op_Explicit(Posit32).0.b_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\;
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := \Quire Posit32::op_Explicit(Posit32).0.return_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.86\ := signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\), 32)) + to_signed(2, 32);
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.87\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.86\ <= to_signed(32, 32);

                        
                        
                        

                        if (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.87\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_67\;
                        else 
                            
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_66\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_64\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.81\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.80\ = \Quire Posit32::op_Explicit(Posit32).0.num_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\;
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.82\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.79\ and \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.81\;
                        if (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.82\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.83\ := shift_left(\Quire Posit32::op_Explicit(Posit32).0.bits_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\, to_integer(unsigned(SmartResize(to_signed(1, 32), 5))));
                            \Quire Posit32::op_Explicit(Posit32).0.bits_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.83\;
                            
                            
                            
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_65\;
                        else 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_63\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_65\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.84\ := SmartResize(unsigned(signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.b_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\), 32)) + to_signed(1, 32)), 8);
                        \Quire Posit32::op_Explicit(Posit32).0.b_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.84\);
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.85\ := \Quire Posit32::op_Explicit(Posit32).0.num2_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ + to_signed(1, 32);
                        \Quire Posit32::op_Explicit(Posit32).0.num2_f9d1c0948957a79ca7758767cdb551a2fd521596e0a020604db70bc0313c407b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.85\;
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_65\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_62\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_66\ => 
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.93\ := to_signed(32, 32) - signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\), 32));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.94\ := SmartResize(unsigned(\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.93\ - to_signed(1, 32)), 8);
                        \Quire Posit32::op_Explicit(Posit32).0.return_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.94\);
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_3\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_67\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.88\ := signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\), 32)) + to_signed(2, 32);
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.89\ := to_signed(32, 32) - (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.88\);
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_68\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_68\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.90\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.89\ > to_signed(2, 32);

                        
                        
                        
                        

                        if ((\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.90\)) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_70\;
                        else 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_71\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_69\ => 
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.return_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := SmartResize(unsigned((\Quire Posit32::op_Explicit(Posit32).0.conditional68bcd4673000ed90d5e5bddf9742548ff8843dd36c272b449a1de261af0ae5a9_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\)), 8);
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_3\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_70\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditional68bcd4673000ed90d5e5bddf9742548ff8843dd36c272b449a1de261af0ae5a9_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := to_signed(2, 32);
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_70\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_69\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_71\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.91\ := signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.b_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\), 32)) + to_signed(2, 32);
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.92\ := SmartResize(unsigned(to_signed(32, 32) - (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.91\)), 8);
                        \Quire Posit32::op_Explicit(Posit32).0.conditional68bcd4673000ed90d5e5bddf9742548ff8843dd36c272b449a1de261af0ae5a9_fa5c7efa4c67d060a70b49e02aabb5ee02fd5c8b1d6e04e5196ceda62f23fe5a\ := signed(SmartResize(((\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.92\)), 32));
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_71\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_69\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_72\ => 
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_72\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_66\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_73\ => 
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.bits_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := (\Quire Posit32::op_Explicit(Posit32).0.conditional963d17004b6788ad55358cce58986fa179ec1b5dc039dfede93d706448099e92_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := \Quire Posit32::op_Explicit(Posit32).0.bits_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\;
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.startingPosition_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := SmartResize(unsigned(to_signed(31, 32)), 8);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.b_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := SmartResize(unsigned(to_signed(1, 32)), 8);
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.98\ := to_signed(32, 32) - signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.startingPosition_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\), 32));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.99\ := shift_left(\Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\, to_integer(unsigned(SmartResize(\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.98\, 5))));
                        \Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.99\;
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_76\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_74\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditional963d17004b6788ad55358cce58986fa179ec1b5dc039dfede93d706448099e92_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := \Quire Posit32::op_Explicit(Posit32).0.this_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\.\PositBits\;
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_74\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_73\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_75\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.bits_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := \Quire Posit32::op_Explicit(Posit32).0.this_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\.\PositBits\;
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.7\ := not(\Quire Posit32::op_Explicit(Posit32).0.bits_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\);
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.97\ := SmartResize(unsigned(signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.unaryOperationResult.7\), 64)) + to_signed(1, 64)), 32);
                        \Quire Posit32::op_Explicit(Posit32).0.return_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.97\);
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditional963d17004b6788ad55358cce58986fa179ec1b5dc039dfede93d706448099e92_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := \Quire Posit32::op_Explicit(Posit32).0.return_c8598ebe73f9f5bfb88d0df855ee308f9c4caf4ef5760e9d645383f544733d31_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\;
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_75\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_73\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_76\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.100\ := shift_right(\Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\, to_integer(unsigned(SmartResize(to_signed(31, 32), 5) and "11111")));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.101\ := (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.100\) and to_unsigned(1, 32);
                        \Quire Posit32::op_Explicit(Posit32).0.num_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.101\;
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.102\ := shift_left(\Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\, to_integer(unsigned(SmartResize(to_signed(1, 32), 5))));
                        \Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.102\;
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.num2_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := to_signed(0, 32);
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_77\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_77\ => 
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.103\ := (\Quire Posit32::op_Explicit(Posit32).0.num2_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\) < signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.startingPosition_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\), 32));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.104\ := shift_right(\Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\, to_integer(unsigned(SmartResize(to_signed(31, 32), 5) and "11111")));
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_79\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_78\ => 
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.return_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := \Quire Posit32::op_Explicit(Posit32).0.b_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\;
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.110\ := signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.return_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\), 32)) + to_signed(2, 32);
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.111\ := SmartResize(\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.110\ + to_signed(2, 32), 32);
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_81\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_79\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.105\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.104\ = \Quire Posit32::op_Explicit(Posit32).0.num_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\;
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.106\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.103\ and \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.105\;
                        if (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.106\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.107\ := shift_left(\Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\, to_integer(unsigned(SmartResize(to_signed(1, 32), 5))));
                            \Quire Posit32::op_Explicit(Posit32).0.bits_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.107\;
                            
                            
                            
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_80\;
                        else 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_78\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_80\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.108\ := SmartResize(unsigned(signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.b_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\), 32)) + to_signed(1, 32)), 8);
                        \Quire Posit32::op_Explicit(Posit32).0.b_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.108\);
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.109\ := \Quire Posit32::op_Explicit(Posit32).0.num2_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ + to_signed(1, 32);
                        \Quire Posit32::op_Explicit(Posit32).0.num2_aa1887a732f44ab7933da762327f79580f968b608eddfcba10dec20b0026fde4_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.109\;
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_80\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_77\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_81\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.112\ := to_signed(32, 32) - (\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.111\);
                        \Quire Posit32::op_Explicit(Posit32).0.num_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.112\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.113\ := \Quire Posit32::op_Explicit(Posit32).0.num_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ > to_signed(0, 32);

                        
                        
                        
                        

                        if ((\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.113\)) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_83\;
                        else 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_84\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_82\ => 
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.return_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := \Quire Posit32::op_Explicit(Posit32).0.conditionalf2eba7c459dd057c9270f346c2a9013399b4309fc21683746ef1be47061f03f1_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\;
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.114\ := shift_right(\Quire Posit32::op_Explicit(Posit32).0.num_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\, to_integer(unsigned(SmartResize(signed(\Quire Posit32::op_Explicit(Posit32).0.return_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\), 5) and "11111")));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.115\ := to_signed(32, 32) - signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.b_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\), 32));
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_85\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_83\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditionalf2eba7c459dd057c9270f346c2a9013399b4309fc21683746ef1be47061f03f1_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := (unsigned(\Quire Posit32::op_Explicit(Posit32).0.num_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\));
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_83\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_82\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_84\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditionalf2eba7c459dd057c9270f346c2a9013399b4309fc21683746ef1be47061f03f1_94bef725a1b90b0f1b2e9d5058b7a34e74ecdb8cab8ec5897a685559b4937cd4\ := to_unsigned(0, 32);
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_84\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_82\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_85\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.116\ := shift_left(\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.114\, to_integer(unsigned(SmartResize(\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.115\, 5))));
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.117\ := shift_right(\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.116\, to_integer(unsigned(SmartResize(to_signed(30, 32), 5) and "11111")));
                        \Quire Posit32::op_Explicit(Posit32).0.num_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.117\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_86\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_86\ => 
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.118\ := signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.b_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\), 32)) /= to_signed(0, 32);

                        
                        
                        
                        

                        if ((\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.118\)) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_88\;
                        else 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_89\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_87\ => 
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.return_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.conditionala233560fe7dfff22c231bec46671f442fee11494dc774056e64d669ec36cdb00_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\;
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.119\ := SmartResize(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.regimeKValue_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\), 32) * to_signed(4, 32), 64);
                        \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.120\ := SmartResize((\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.119\) + signed(SmartResize((\Quire Posit32::op_Explicit(Posit32).0.return_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\), 64)), 16);
                        \Quire Posit32::op_Explicit(Posit32).0.conditional1aa95b35288eb627929161a1ee637479589960934567100c958634e64afb13de_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := SmartResize(((\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.120\)), 32);
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_87\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_53\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_88\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditionala233560fe7dfff22c231bec46671f442fee11494dc774056e64d669ec36cdb00_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := \Quire Posit32::op_Explicit(Posit32).0.num_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\;
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_88\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_87\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_89\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditionala233560fe7dfff22c231bec46671f442fee11494dc774056e64d669ec36cdb00_b30c7cf04e18e8e1d9326fda65a98f3e6ce2cb9a087dd14bb74739b64c0a2a6c_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_unsigned(0, 32);
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_89\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_87\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_90\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.conditional1aa95b35288eb627929161a1ee637479589960934567100c958634e64afb13de_5547e2b2a08e312134cbdc7a0930a7319e6155fa1d1d0c7cedcf0662fda61e28\ := to_signed(0, 32);
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_90\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_53\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_91\ => 
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ = \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\) then 
                            \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ <= false;
                            \Quire Posit32::op_Explicit(Posit32).0.return.1\ := \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).return.0\;
                            \Quire Posit32::op_Explicit(Posit32).0.quire\ := \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.In.0\;
                            \Quire Posit32::op_Explicit(Posit32).0.quire\ := \Quire Posit32::op_Explicit(Posit32).0.return.1\;
                            
                            
                            
                            
                            
                            
                            \Quire Posit32::op_Explicit(Posit32).0.this_5204dd194817ce0e22c54ac6e6fe7dc0a0e40352e5a5fed887c54294684dded0\ := \Quire Posit32::op_Explicit(Posit32).0.x\;
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.123\ := signed(SmartResize(\Quire Posit32::op_Explicit(Posit32).0.this_5204dd194817ce0e22c54ac6e6fe7dc0a0e40352e5a5fed887c54294684dded0\.\PositBits\ and "10000000000000000000000000000000", 64));
                            \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.124\ := signed(SmartResize(((\Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.123\)), 64)) = to_signed(0, 64);
                            \Quire Posit32::op_Explicit(Posit32).0.return_5204dd194817ce0e22c54ac6e6fe7dc0a0e40352e5a5fed887c54294684dded0\ := \Quire Posit32::op_Explicit(Posit32).0.binaryOperationResult.124\;
                            
                            
                            
                            
                            

                            
                            
                            

                            if (\Quire Posit32::op_Explicit(Posit32).0.return_5204dd194817ce0e22c54ac6e6fe7dc0a0e40352e5a5fed887c54294684dded0\) then 
                                \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_93\;
                            else 
                                
                                \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_92\;
                            end if;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_92\ => 
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_OnesComplement(Quire).q.parameter.Out.0\ <= \Quire Posit32::op_Explicit(Posit32).0.quire\;
                        \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_OnesComplement(Quire)._Started.0\ <= true;
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_94\;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_93\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Posit32::op_Explicit(Posit32).0.return\ <= \Quire Posit32::op_Explicit(Posit32).0.quire\;
                        \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_1\;
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0._State\ = \Quire Posit32::op_Explicit(Posit32).0._State_93\) then 
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_92\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_94\ => 
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_OnesComplement(Quire)._Started.0\ = \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_OnesComplement(Quire)._Finished.0\) then 
                            \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_OnesComplement(Quire)._Started.0\ <= false;
                            \Quire Posit32::op_Explicit(Posit32).0.return.2\ := \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_OnesComplement(Quire).return.0\;
                            \Quire Posit32::op_Explicit(Posit32).0.quire\ := \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_OnesComplement(Quire).q.parameter.In.0\;
                            
                            \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32).left.parameter.Out.0\ <= \Quire Posit32::op_Explicit(Posit32).0.return.2\;
                            \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32).right.parameter.Out.0\ <= to_unsigned(1, 32);
                            \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32)._Started.0\ <= true;
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_95\;
                        end if;
                        
                    when \Quire Posit32::op_Explicit(Posit32).0._State_95\ => 
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32)._Started.0\ = \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32)._Finished.0\) then 
                            \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32)._Started.0\ <= false;
                            \Quire Posit32::op_Explicit(Posit32).0.return.3\ := \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32).return.0\;
                            \Quire Posit32::op_Explicit(Posit32).0.return.2\ := \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32).left.parameter.In.0\;
                            \Quire Posit32::op_Explicit(Posit32).0.return\ <= \Quire Posit32::op_Explicit(Posit32).0.return.3\;
                            \Quire Posit32::op_Explicit(Posit32).0._State\ := \Quire Posit32::op_Explicit(Posit32).0._State_1\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Quire::.ctor(UInt64[],UInt16).0._StateMachine\: process (\Clock\) 
        Variable \Quire::.ctor(UInt64[],UInt16).0._State\: \Quire::.ctor(UInt64[],UInt16).0._States\ := \Quire::.ctor(UInt64[],UInt16).0._State_0\;
        Variable \Quire::.ctor(UInt64[],UInt16).0.this\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire::.ctor(UInt64[],UInt16).0.segments\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
        Variable \Quire::.ctor(UInt64[],UInt16).0.size\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire::.ctor(UInt64[],UInt16).0.num\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire::.ctor(UInt64[],UInt16).0.binaryOperationResult.0\: boolean := false;
        Variable \Quire::.ctor(UInt64[],UInt16).0.binaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Quire::.ctor(UInt64[],UInt16).0._Finished\ <= false;
                \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.Out\ <= (others => to_unsigned(0, 64));
                \Quire::.ctor(UInt64[],UInt16).0._State\ := \Quire::.ctor(UInt64[],UInt16).0._State_0\;
                \Quire::.ctor(UInt64[],UInt16).0.segments\ := (others => to_unsigned(0, 64));
                \Quire::.ctor(UInt64[],UInt16).0.size\ := to_unsigned(0, 16);
                \Quire::.ctor(UInt64[],UInt16).0.num\ := to_signed(0, 32);
                \Quire::.ctor(UInt64[],UInt16).0.binaryOperationResult.0\ := false;
                \Quire::.ctor(UInt64[],UInt16).0.binaryOperationResult.1\ := to_signed(0, 32);
            else 
                case \Quire::.ctor(UInt64[],UInt16).0._State\ is 
                    when \Quire::.ctor(UInt64[],UInt16).0._State_0\ => 
                        
                        
                        if (\Quire::.ctor(UInt64[],UInt16).0._Started\ = true) then 
                            \Quire::.ctor(UInt64[],UInt16).0._State\ := \Quire::.ctor(UInt64[],UInt16).0._State_2\;
                        end if;
                        
                    when \Quire::.ctor(UInt64[],UInt16).0._State_1\ => 
                        
                        
                        if (\Quire::.ctor(UInt64[],UInt16).0._Started\ = true) then 
                            \Quire::.ctor(UInt64[],UInt16).0._Finished\ <= true;
                        else 
                            \Quire::.ctor(UInt64[],UInt16).0._Finished\ <= false;
                            \Quire::.ctor(UInt64[],UInt16).0._State\ := \Quire::.ctor(UInt64[],UInt16).0._State_0\;
                        end if;
                        
                        \Quire::.ctor(UInt64[],UInt16).0.this.parameter.Out\ <= \Quire::.ctor(UInt64[],UInt16).0.this\;
                        \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.Out\ <= \Quire::.ctor(UInt64[],UInt16).0.segments\;
                        
                    when \Quire::.ctor(UInt64[],UInt16).0._State_2\ => 
                        \Quire::.ctor(UInt64[],UInt16).0.this\ := \Quire::.ctor(UInt64[],UInt16).0.this.parameter.In\;
                        \Quire::.ctor(UInt64[],UInt16).0.segments\ := \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.In\;
                        \Quire::.ctor(UInt64[],UInt16).0.size\ := \Quire::.ctor(UInt64[],UInt16).0.size.parameter.In\;
                        
                        
                        
                        \Quire::.ctor(UInt64[],UInt16).0.this\.\SegmentCount\ := to_unsigned(8, 16);
                        
                        
                        
                        \Quire::.ctor(UInt64[],UInt16).0.this\.\Size\ := SmartResize(unsigned(to_signed(0, 32)), 16);
                        
                        
                        
                        \Quire::.ctor(UInt64[],UInt16).0.this\.\Segments\ := (others => to_unsigned(0, 64));
                        
                        
                        
                        \Quire::.ctor(UInt64[],UInt16).0.this\.\Segments\ := \Quire::.ctor(UInt64[],UInt16).0.segments\(0 to 7);
                        
                        
                        
                        
                        
                        
                        \Quire::.ctor(UInt64[],UInt16).0.num\ := to_signed(8, 32);
                        
                        
                        
                        
                        
                        
                        
                        \Quire::.ctor(UInt64[],UInt16).0._State\ := \Quire::.ctor(UInt64[],UInt16).0._State_3\;
                        
                    when \Quire::.ctor(UInt64[],UInt16).0._State_3\ => 
                        
                        
                        \Quire::.ctor(UInt64[],UInt16).0.binaryOperationResult.0\ := (\Quire::.ctor(UInt64[],UInt16).0.num\) < to_signed(8, 32);
                        if (\Quire::.ctor(UInt64[],UInt16).0.binaryOperationResult.0\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire::.ctor(UInt64[],UInt16).0.this\.\Segments\(to_integer(\Quire::.ctor(UInt64[],UInt16).0.num\)) := to_unsigned(0, 64);
                            
                            
                            
                            \Quire::.ctor(UInt64[],UInt16).0.binaryOperationResult.1\ := \Quire::.ctor(UInt64[],UInt16).0.num\ + to_signed(1, 32);
                            \Quire::.ctor(UInt64[],UInt16).0.num\ := \Quire::.ctor(UInt64[],UInt16).0.binaryOperationResult.1\;
                        else 
                            \Quire::.ctor(UInt64[],UInt16).0._State\ := \Quire::.ctor(UInt64[],UInt16).0._State_4\;
                        end if;
                        
                    when \Quire::.ctor(UInt64[],UInt16).0._State_4\ => 
                        
                        \Quire::.ctor(UInt64[],UInt16).0._State\ := \Quire::.ctor(UInt64[],UInt16).0._State_1\;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Quire::.ctor(UInt32,UInt16).0._StateMachine\: process (\Clock\) 
        Variable \Quire::.ctor(UInt32,UInt16).0._State\: \Quire::.ctor(UInt32,UInt16).0._States\ := \Quire::.ctor(UInt32,UInt16).0._State_0\;
        Variable \Quire::.ctor(UInt32,UInt16).0.this\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire::.ctor(UInt32,UInt16).0.firstSegment\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire::.ctor(UInt32,UInt16).0.size\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire::.ctor(UInt32,UInt16).0.conditional508ca86de85a5da84bb49b246fc4b145e1352a0547a47e41f17ab54c68695517\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire::.ctor(UInt32,UInt16).0.remainderOperand0c439d9dfdc1e321f9179f8d0530a346aae5aa4d433af564a6e961f787b90b5b\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.3\: boolean := false;
        Variable \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.4\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.5\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire::.ctor(UInt32,UInt16).0.num\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.6\: boolean := false;
        Variable \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.7\: signed(31 downto 0) := to_signed(0, 32);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Quire::.ctor(UInt32,UInt16).0._Finished\ <= false;
                \Quire::.ctor(UInt32,UInt16).0._State\ := \Quire::.ctor(UInt32,UInt16).0._State_0\;
                \Quire::.ctor(UInt32,UInt16).0.firstSegment\ := to_unsigned(0, 32);
                \Quire::.ctor(UInt32,UInt16).0.size\ := to_unsigned(0, 16);
                \Quire::.ctor(UInt32,UInt16).0.conditional508ca86de85a5da84bb49b246fc4b145e1352a0547a47e41f17ab54c68695517\ := to_signed(0, 32);
                \Quire::.ctor(UInt32,UInt16).0.remainderOperand0c439d9dfdc1e321f9179f8d0530a346aae5aa4d433af564a6e961f787b90b5b\ := to_signed(0, 32);
                \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.0\ := to_signed(0, 32);
                \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.1\ := to_signed(0, 32);
                \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.2\ := to_signed(0, 32);
                \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.3\ := false;
                \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.4\ := to_signed(0, 32);
                \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.5\ := to_unsigned(0, 16);
                \Quire::.ctor(UInt32,UInt16).0.num\ := to_signed(0, 32);
                \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.6\ := false;
                \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.7\ := to_signed(0, 32);
            else 
                case \Quire::.ctor(UInt32,UInt16).0._State\ is 
                    when \Quire::.ctor(UInt32,UInt16).0._State_0\ => 
                        
                        
                        if (\Quire::.ctor(UInt32,UInt16).0._Started\ = true) then 
                            \Quire::.ctor(UInt32,UInt16).0._State\ := \Quire::.ctor(UInt32,UInt16).0._State_2\;
                        end if;
                        
                    when \Quire::.ctor(UInt32,UInt16).0._State_1\ => 
                        
                        
                        if (\Quire::.ctor(UInt32,UInt16).0._Started\ = true) then 
                            \Quire::.ctor(UInt32,UInt16).0._Finished\ <= true;
                        else 
                            \Quire::.ctor(UInt32,UInt16).0._Finished\ <= false;
                            \Quire::.ctor(UInt32,UInt16).0._State\ := \Quire::.ctor(UInt32,UInt16).0._State_0\;
                        end if;
                        
                        \Quire::.ctor(UInt32,UInt16).0.this.parameter.Out\ <= \Quire::.ctor(UInt32,UInt16).0.this\;
                        
                    when \Quire::.ctor(UInt32,UInt16).0._State_2\ => 
                        \Quire::.ctor(UInt32,UInt16).0.this\ := \Quire::.ctor(UInt32,UInt16).0.this.parameter.In\;
                        \Quire::.ctor(UInt32,UInt16).0.firstSegment\ := \Quire::.ctor(UInt32,UInt16).0.firstSegment.parameter.In\;
                        \Quire::.ctor(UInt32,UInt16).0.size\ := \Quire::.ctor(UInt32,UInt16).0.size.parameter.In\;
                        
                        
                        
                        \Quire::.ctor(UInt32,UInt16).0.this\.\Size\ := \Quire::.ctor(UInt32,UInt16).0.size\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire::.ctor(UInt32,UInt16).0.remainderOperand0c439d9dfdc1e321f9179f8d0530a346aae5aa4d433af564a6e961f787b90b5b\ := signed(SmartResize(\Quire::.ctor(UInt32,UInt16).0.size\, 32));
                        
                        
                        
                        
                        
                        
                        
                        \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.0\ := \Quire::.ctor(UInt32,UInt16).0.remainderOperand0c439d9dfdc1e321f9179f8d0530a346aae5aa4d433af564a6e961f787b90b5b\ / to_signed(32, 32);
                        \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.1\ := SmartResize(\Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.0\ * to_signed(32, 32), 32);
                        \Quire::.ctor(UInt32,UInt16).0._State\ := \Quire::.ctor(UInt32,UInt16).0._State_3\;
                        
                    when \Quire::.ctor(UInt32,UInt16).0._State_3\ => 
                        
                        \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.2\ := \Quire::.ctor(UInt32,UInt16).0.remainderOperand0c439d9dfdc1e321f9179f8d0530a346aae5aa4d433af564a6e961f787b90b5b\ - \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.1\;
                        \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.3\ := \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.2\ /= to_signed(0, 32);

                        
                        
                        
                        

                        if ((\Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.3\)) then 
                            \Quire::.ctor(UInt32,UInt16).0._State\ := \Quire::.ctor(UInt32,UInt16).0._State_5\;
                        else 
                            \Quire::.ctor(UInt32,UInt16).0._State\ := \Quire::.ctor(UInt32,UInt16).0._State_6\;
                        end if;
                        
                    when \Quire::.ctor(UInt32,UInt16).0._State_4\ => 
                        
                        
                        
                        
                        \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.4\ := shift_right(signed(SmartResize((\Quire::.ctor(UInt32,UInt16).0.size\), 32)), to_integer(unsigned(SmartResize(to_signed(6, 32), 5) and "11111")));
                        \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.5\ := SmartResize(unsigned((\Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.4\) + (\Quire::.ctor(UInt32,UInt16).0.conditional508ca86de85a5da84bb49b246fc4b145e1352a0547a47e41f17ab54c68695517\)), 16);
                        \Quire::.ctor(UInt32,UInt16).0.this\.\SegmentCount\ := (\Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.5\);
                        
                        
                        
                        \Quire::.ctor(UInt32,UInt16).0.this\.\Segments\ := (others => to_unsigned(0, 64));
                        
                        
                        
                        \Quire::.ctor(UInt32,UInt16).0.this\.\Segments\(to_integer(to_signed(0, 32))) := SmartResize(to_unsigned(1, 32), 64);
                        
                        
                        
                        
                        
                        
                        \Quire::.ctor(UInt32,UInt16).0.num\ := to_signed(1, 32);
                        
                        
                        
                        
                        
                        
                        
                        \Quire::.ctor(UInt32,UInt16).0._State\ := \Quire::.ctor(UInt32,UInt16).0._State_7\;
                        
                    when \Quire::.ctor(UInt32,UInt16).0._State_5\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire::.ctor(UInt32,UInt16).0.conditional508ca86de85a5da84bb49b246fc4b145e1352a0547a47e41f17ab54c68695517\ := to_signed(1, 32);
                        
                        if (\Quire::.ctor(UInt32,UInt16).0._State\ = \Quire::.ctor(UInt32,UInt16).0._State_5\) then 
                            \Quire::.ctor(UInt32,UInt16).0._State\ := \Quire::.ctor(UInt32,UInt16).0._State_4\;
                        end if;
                        
                    when \Quire::.ctor(UInt32,UInt16).0._State_6\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire::.ctor(UInt32,UInt16).0.conditional508ca86de85a5da84bb49b246fc4b145e1352a0547a47e41f17ab54c68695517\ := to_signed(0, 32);
                        
                        if (\Quire::.ctor(UInt32,UInt16).0._State\ = \Quire::.ctor(UInt32,UInt16).0._State_6\) then 
                            \Quire::.ctor(UInt32,UInt16).0._State\ := \Quire::.ctor(UInt32,UInt16).0._State_4\;
                        end if;
                        
                    when \Quire::.ctor(UInt32,UInt16).0._State_7\ => 
                        
                        
                        \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.6\ := (\Quire::.ctor(UInt32,UInt16).0.num\) < signed(SmartResize((\Quire::.ctor(UInt32,UInt16).0.this\.\SegmentCount\), 32));
                        if (\Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.6\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire::.ctor(UInt32,UInt16).0.this\.\Segments\(to_integer(\Quire::.ctor(UInt32,UInt16).0.num\)) := to_unsigned(0, 64);
                            
                            
                            
                            \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.7\ := \Quire::.ctor(UInt32,UInt16).0.num\ + to_signed(1, 32);
                            \Quire::.ctor(UInt32,UInt16).0.num\ := \Quire::.ctor(UInt32,UInt16).0.binaryOperationResult.7\;
                        else 
                            \Quire::.ctor(UInt32,UInt16).0._State\ := \Quire::.ctor(UInt32,UInt16).0._State_8\;
                        end if;
                        
                    when \Quire::.ctor(UInt32,UInt16).0._State_8\ => 
                        
                        \Quire::.ctor(UInt32,UInt16).0._State\ := \Quire::.ctor(UInt32,UInt16).0._State_1\;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Quire Quire::op_Addition(Quire,Quire).0._StateMachine\: process (\Clock\) 
        Variable \Quire Quire::op_Addition(Quire,Quire).0._State\: \Quire Quire::op_Addition(Quire,Quire).0._States\ := \Quire Quire::op_Addition(Quire,Quire).0._State_0\;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.left\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.right\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.0\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.1\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.2\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.array\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
        Variable \Quire Quire::op_Addition(Quire,Quire).0.flag\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.num\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.num2\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.num3\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.3\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.4\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.flag2\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.5\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.6\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.7\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.flag3\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.8\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.9\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.10\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.b\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.conditional746a1c636f616ff3623be4e48942688719382078a087cbdab0e2c998303da9ba\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.conditionalc042a0f1121d35344a49419953dc5f52591ee75c13d7b4714794eeff7d14bf49\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.conditionalae2b32de30beca2038d02dc985eb3cd14f87df2ffaa1520711b83d6b5e0acd70\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.11\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.12\: unsigned(7 downto 0) := to_unsigned(0, 8);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.13\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.14\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.15\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.16\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.17\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.18\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.19\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.20\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.21\: boolean := false;
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.22\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.23\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_Addition(Quire,Quire).0.objectd7f66d6090a3f51dbf9c6b85d3744cbaf909687ec9d3f52027672e9a5e2ece9d\: \Lombiq.Arithmetics.Quire\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Quire Quire::op_Addition(Quire,Quire).0._Finished\ <= false;
                \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 64));
                \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= false;
                \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_0\;
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.0\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.1\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.2\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.array\ := (others => to_unsigned(0, 64));
                \Quire Quire::op_Addition(Quire,Quire).0.flag\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.num\ := to_unsigned(0, 16);
                \Quire Quire::op_Addition(Quire,Quire).0.num2\ := to_unsigned(0, 16);
                \Quire Quire::op_Addition(Quire,Quire).0.num3\ := to_unsigned(0, 16);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.3\ := to_signed(0, 32);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.4\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.flag2\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.5\ := to_unsigned(0, 64);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.6\ := to_unsigned(0, 64);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.7\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.flag3\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.8\ := to_unsigned(0, 64);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.9\ := to_unsigned(0, 64);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.10\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.b\ := to_unsigned(0, 8);
                \Quire Quire::op_Addition(Quire,Quire).0.conditional746a1c636f616ff3623be4e48942688719382078a087cbdab0e2c998303da9ba\ := to_signed(0, 32);
                \Quire Quire::op_Addition(Quire,Quire).0.conditionalc042a0f1121d35344a49419953dc5f52591ee75c13d7b4714794eeff7d14bf49\ := to_signed(0, 32);
                \Quire Quire::op_Addition(Quire,Quire).0.conditionalae2b32de30beca2038d02dc985eb3cd14f87df2ffaa1520711b83d6b5e0acd70\ := to_signed(0, 32);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.11\ := to_signed(0, 32);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.12\ := to_unsigned(0, 8);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.13\ := to_signed(0, 32);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.14\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.15\ := to_unsigned(0, 64);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.16\ := to_unsigned(0, 64);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.17\ := to_signed(0, 32);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.18\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.19\ := to_unsigned(0, 16);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.20\ := to_signed(0, 32);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.21\ := false;
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.22\ := to_unsigned(0, 16);
                \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.23\ := to_unsigned(0, 16);
            else 
                case \Quire Quire::op_Addition(Quire,Quire).0._State\ is 
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_0\ => 
                        
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._Started\ = true) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_2\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_1\ => 
                        
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._Started\ = true) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._Finished\ <= true;
                        else 
                            \Quire Quire::op_Addition(Quire,Quire).0._Finished\ <= false;
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_0\;
                        end if;
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.left.parameter.Out\ <= \Quire Quire::op_Addition(Quire,Quire).0.left\;
                        \Quire Quire::op_Addition(Quire,Quire).0.right.parameter.Out\ <= \Quire Quire::op_Addition(Quire,Quire).0.right\;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_2\ => 
                        \Quire Quire::op_Addition(Quire,Quire).0.left\ := \Quire Quire::op_Addition(Quire,Quire).0.left.parameter.In\;
                        \Quire Quire::op_Addition(Quire,Quire).0.right\ := \Quire Quire::op_Addition(Quire,Quire).0.right.parameter.In\;
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.0\ := signed(SmartResize((\Quire Quire::op_Addition(Quire,Quire).0.left\.\SegmentCount\), 32)) = to_signed(0, 32);
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.1\ := signed(SmartResize((\Quire Quire::op_Addition(Quire,Quire).0.right\.\SegmentCount\), 32)) = to_signed(0, 32);
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.2\ := \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.0\ or \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.1\;

                        
                        
                        

                        if (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.2\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_4\;
                        else 
                            
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_3\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_3\ => 
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.array\ := (others => to_unsigned(0, 64));
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.flag\ := false;
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.num\ := SmartResize(unsigned(to_signed(0, 32)), 16);
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.num2\ := SmartResize(unsigned(to_signed(0, 32)), 16);
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.num3\ := SmartResize(unsigned(to_signed(0, 32)), 16);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_5\;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_4\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.return\ <= \Quire Quire::op_Addition(Quire,Quire).0.left\;
                        \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_1\;
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._State\ = \Quire Quire::op_Addition(Quire,Quire).0._State_4\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_3\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_5\ => 
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.3\ := shift_left(signed(SmartResize((\Quire Quire::op_Addition(Quire,Quire).0.left\.\SegmentCount\), 32)), to_integer(unsigned(SmartResize(to_signed(6, 32), 5))));
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.4\ := signed(SmartResize((\Quire Quire::op_Addition(Quire,Quire).0.num3\), 32)) < (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.3\);
                        if (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.4\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_7\;
                        else 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_6\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_6\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.objectd7f66d6090a3f51dbf9c6b85d3744cbaf909687ec9d3f52027672e9a5e2ece9d\.\IsNull\ := false;
                        \Quire Quire::op_Addition(Quire,Quire).0.objectd7f66d6090a3f51dbf9c6b85d3744cbaf909687ec9d3f52027672e9a5e2ece9d\.\Size\ := to_unsigned(0, 16);
                        \Quire Quire::op_Addition(Quire,Quire).0.objectd7f66d6090a3f51dbf9c6b85d3744cbaf909687ec9d3f52027672e9a5e2ece9d\.\SegmentCount\ := to_unsigned(0, 16);
                        \Quire Quire::op_Addition(Quire,Quire).0.objectd7f66d6090a3f51dbf9c6b85d3744cbaf909687ec9d3f52027672e9a5e2ece9d\.\Segments\ := (others => to_unsigned(0, 64));
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\ <= \Quire Quire::op_Addition(Quire,Quire).0.objectd7f66d6090a3f51dbf9c6b85d3744cbaf909687ec9d3f52027672e9a5e2ece9d\;
                        \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\ <= \Quire Quire::op_Addition(Quire,Quire).0.array\;
                        \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\ <= SmartResize(unsigned(to_signed(0, 32)), 16);
                        \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= true;
                        \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_28\;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_7\ => 
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.5\ := SmartResize(shift_right(\Quire Quire::op_Addition(Quire,Quire).0.left\.\Segments\(to_integer(\Quire Quire::op_Addition(Quire,Quire).0.num\)), to_integer(unsigned(SmartResize(signed(SmartResize(\Quire Quire::op_Addition(Quire,Quire).0.num2\, 32)), 6) and "111111"))), 64);
                        \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_8\;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_8\ => 
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.6\ := (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.5\) and to_unsigned(1, 64);
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.7\ := (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.6\) = to_unsigned(1, 64);
                        \Quire Quire::op_Addition(Quire,Quire).0.flag2\ := \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.7\;
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_9\;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_9\ => 
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.8\ := SmartResize(shift_right(\Quire Quire::op_Addition(Quire,Quire).0.right\.\Segments\(to_integer(\Quire Quire::op_Addition(Quire,Quire).0.num\)), to_integer(unsigned(SmartResize(signed(SmartResize(\Quire Quire::op_Addition(Quire,Quire).0.num2\, 32)), 6) and "111111"))), 64);
                        \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_10\;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_10\ => 
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.9\ := (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.8\) and to_unsigned(1, 64);
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.10\ := (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.9\) = to_unsigned(1, 64);
                        \Quire Quire::op_Addition(Quire,Quire).0.flag3\ := \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.10\;
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        

                        
                        
                        
                        

                        if (\Quire Quire::op_Addition(Quire,Quire).0.flag2\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_12\;
                        else 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_13\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_11\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        

                        
                        
                        
                        

                        if (\Quire Quire::op_Addition(Quire,Quire).0.flag3\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_15\;
                        else 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_16\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_12\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.conditional746a1c636f616ff3623be4e48942688719382078a087cbdab0e2c998303da9ba\ := to_signed(1, 32);
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._State\ = \Quire Quire::op_Addition(Quire,Quire).0._State_12\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_11\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_13\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.conditional746a1c636f616ff3623be4e48942688719382078a087cbdab0e2c998303da9ba\ := to_signed(0, 32);
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._State\ = \Quire Quire::op_Addition(Quire,Quire).0._State_13\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_11\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_14\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        

                        
                        
                        
                        

                        if (\Quire Quire::op_Addition(Quire,Quire).0.flag\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_18\;
                        else 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_19\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_15\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.conditionalc042a0f1121d35344a49419953dc5f52591ee75c13d7b4714794eeff7d14bf49\ := to_signed(1, 32);
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._State\ = \Quire Quire::op_Addition(Quire,Quire).0._State_15\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_14\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_16\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.conditionalc042a0f1121d35344a49419953dc5f52591ee75c13d7b4714794eeff7d14bf49\ := to_signed(0, 32);
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._State\ = \Quire Quire::op_Addition(Quire,Quire).0._State_16\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_14\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_17\ => 
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.11\ := (\Quire Quire::op_Addition(Quire,Quire).0.conditional746a1c636f616ff3623be4e48942688719382078a087cbdab0e2c998303da9ba\) + (\Quire Quire::op_Addition(Quire,Quire).0.conditionalc042a0f1121d35344a49419953dc5f52591ee75c13d7b4714794eeff7d14bf49\);
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.12\ := SmartResize(unsigned(\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.11\ + (\Quire Quire::op_Addition(Quire,Quire).0.conditionalae2b32de30beca2038d02dc985eb3cd14f87df2ffaa1520711b83d6b5e0acd70\)), 8);
                        \Quire Quire::op_Addition(Quire,Quire).0.b\ := (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.12\);
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.13\ := signed(SmartResize((\Quire Quire::op_Addition(Quire,Quire).0.b\), 32)) and to_signed(1, 32);
                        \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_20\;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_18\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.conditionalae2b32de30beca2038d02dc985eb3cd14f87df2ffaa1520711b83d6b5e0acd70\ := to_signed(1, 32);
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._State\ = \Quire Quire::op_Addition(Quire,Quire).0._State_18\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_17\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_19\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.conditionalae2b32de30beca2038d02dc985eb3cd14f87df2ffaa1520711b83d6b5e0acd70\ := to_signed(0, 32);
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._State\ = \Quire Quire::op_Addition(Quire,Quire).0._State_19\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_17\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_20\ => 
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.14\ := (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.13\) = to_signed(1, 32);

                        
                        
                        

                        if (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.14\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_22\;
                        else 
                            
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_21\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_21\ => 
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.17\ := shift_right(signed(SmartResize((\Quire Quire::op_Addition(Quire,Quire).0.b\), 32)), to_integer(unsigned(SmartResize(to_signed(1, 32), 5) and "11111")));
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.18\ := \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.17\ = to_signed(1, 32);
                        \Quire Quire::op_Addition(Quire,Quire).0.flag\ := \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.18\;
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_24\;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_22\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.15\ := SmartResize(unsigned(shift_left(to_signed(1, 64), to_integer(unsigned(SmartResize(signed(SmartResize(\Quire Quire::op_Addition(Quire,Quire).0.num2\, 32)), 6))))), 64);
                        \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_23\;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_23\ => 
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.16\ := \Quire Quire::op_Addition(Quire,Quire).0.array\(to_integer(\Quire Quire::op_Addition(Quire,Quire).0.num\)) + (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.15\);
                        \Quire Quire::op_Addition(Quire,Quire).0.array\(to_integer(\Quire Quire::op_Addition(Quire,Quire).0.num\)) := \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.16\;
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._State\ = \Quire Quire::op_Addition(Quire,Quire).0._State_23\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_21\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_24\ => 
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.19\ := SmartResize(unsigned(signed(SmartResize((\Quire Quire::op_Addition(Quire,Quire).0.num2\), 32)) + to_signed(1, 32)), 16);
                        \Quire Quire::op_Addition(Quire,Quire).0.num2\ := (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.19\);
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.20\ := shift_right(signed(SmartResize((\Quire Quire::op_Addition(Quire,Quire).0.num2\), 32)), to_integer(unsigned(SmartResize(to_signed(6, 32), 5) and "11111")));
                        \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_25\;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_25\ => 
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.21\ := \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.20\ = to_signed(1, 32);

                        
                        
                        

                        if (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.21\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_27\;
                        else 
                            
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_26\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_26\ => 
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.23\ := SmartResize(unsigned(signed(SmartResize((\Quire Quire::op_Addition(Quire,Quire).0.num3\), 32)) + to_signed(1, 32)), 16);
                        \Quire Quire::op_Addition(Quire,Quire).0.num3\ := (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.23\);
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._State\ = \Quire Quire::op_Addition(Quire,Quire).0._State_26\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_5\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_27\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.num2\ := SmartResize(unsigned(to_signed(0, 32)), 16);
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.22\ := SmartResize(unsigned(signed(SmartResize((\Quire Quire::op_Addition(Quire,Quire).0.num\), 32)) + to_signed(1, 32)), 16);
                        \Quire Quire::op_Addition(Quire,Quire).0.num\ := (\Quire Quire::op_Addition(Quire,Quire).0.binaryOperationResult.22\);
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0._State\ = \Quire Quire::op_Addition(Quire,Quire).0._State_27\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_26\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,Quire).0._State_28\ => 
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ = \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= false;
                            \Quire Quire::op_Addition(Quire,Quire).0.objectd7f66d6090a3f51dbf9c6b85d3744cbaf909687ec9d3f52027672e9a5e2ece9d\ := \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\;
                            \Quire Quire::op_Addition(Quire,Quire).0.array\ := \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\;
                            
                            
                            
                            \Quire Quire::op_Addition(Quire,Quire).0.return\ <= \Quire Quire::op_Addition(Quire,Quire).0.objectd7f66d6090a3f51dbf9c6b85d3744cbaf909687ec9d3f52027672e9a5e2ece9d\;
                            \Quire Quire::op_Addition(Quire,Quire).0._State\ := \Quire Quire::op_Addition(Quire,Quire).0._State_1\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Quire Quire::op_Addition(Quire,UInt32).0._StateMachine\: process (\Clock\) 
        Variable \Quire Quire::op_Addition(Quire,UInt32).0._State\: \Quire Quire::op_Addition(Quire,UInt32).0._States\ := \Quire Quire::op_Addition(Quire,UInt32).0._State_0\;
        Variable \Quire Quire::op_Addition(Quire,UInt32).0.left\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire Quire::op_Addition(Quire,UInt32).0.right\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Quire::op_Addition(Quire,UInt32).0.object2b25f3fa9b50e7492d78b34e15a583b8300db89f75b5c7cb2910bbab85a19ff0\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire Quire::op_Addition(Quire,UInt32).0.binaryOperationResult.0\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_Addition(Quire,UInt32).0.return.0\: \Lombiq.Arithmetics.Quire\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Quire Quire::op_Addition(Quire,UInt32).0._Finished\ <= false;
                \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).firstSegment.parameter.Out.0\ <= to_unsigned(0, 32);
                \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Started.0\ <= false;
                \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\ <= false;
                \Quire Quire::op_Addition(Quire,UInt32).0._State\ := \Quire Quire::op_Addition(Quire,UInt32).0._State_0\;
                \Quire Quire::op_Addition(Quire,UInt32).0.right\ := to_unsigned(0, 32);
                \Quire Quire::op_Addition(Quire,UInt32).0.binaryOperationResult.0\ := to_unsigned(0, 16);
            else 
                case \Quire Quire::op_Addition(Quire,UInt32).0._State\ is 
                    when \Quire Quire::op_Addition(Quire,UInt32).0._State_0\ => 
                        
                        
                        if (\Quire Quire::op_Addition(Quire,UInt32).0._Started\ = true) then 
                            \Quire Quire::op_Addition(Quire,UInt32).0._State\ := \Quire Quire::op_Addition(Quire,UInt32).0._State_2\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,UInt32).0._State_1\ => 
                        
                        
                        if (\Quire Quire::op_Addition(Quire,UInt32).0._Started\ = true) then 
                            \Quire Quire::op_Addition(Quire,UInt32).0._Finished\ <= true;
                        else 
                            \Quire Quire::op_Addition(Quire,UInt32).0._Finished\ <= false;
                            \Quire Quire::op_Addition(Quire,UInt32).0._State\ := \Quire Quire::op_Addition(Quire,UInt32).0._State_0\;
                        end if;
                        
                        \Quire Quire::op_Addition(Quire,UInt32).0.left.parameter.Out\ <= \Quire Quire::op_Addition(Quire,UInt32).0.left\;
                        
                    when \Quire Quire::op_Addition(Quire,UInt32).0._State_2\ => 
                        \Quire Quire::op_Addition(Quire,UInt32).0.left\ := \Quire Quire::op_Addition(Quire,UInt32).0.left.parameter.In\;
                        \Quire Quire::op_Addition(Quire,UInt32).0.right\ := \Quire Quire::op_Addition(Quire,UInt32).0.right.parameter.In\;
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_Addition(Quire,UInt32).0.object2b25f3fa9b50e7492d78b34e15a583b8300db89f75b5c7cb2910bbab85a19ff0\.\IsNull\ := false;
                        \Quire Quire::op_Addition(Quire,UInt32).0.object2b25f3fa9b50e7492d78b34e15a583b8300db89f75b5c7cb2910bbab85a19ff0\.\Size\ := to_unsigned(0, 16);
                        \Quire Quire::op_Addition(Quire,UInt32).0.object2b25f3fa9b50e7492d78b34e15a583b8300db89f75b5c7cb2910bbab85a19ff0\.\SegmentCount\ := to_unsigned(0, 16);
                        \Quire Quire::op_Addition(Quire,UInt32).0.object2b25f3fa9b50e7492d78b34e15a583b8300db89f75b5c7cb2910bbab85a19ff0\.\Segments\ := (others => to_unsigned(0, 64));
                        
                        \Quire Quire::op_Addition(Quire,UInt32).0.binaryOperationResult.0\ := SmartResize(unsigned(shift_left(signed(SmartResize((\Quire Quire::op_Addition(Quire,UInt32).0.left\.\SegmentCount\), 32)), to_integer(unsigned(SmartResize(to_signed(6, 32), 5))))), 16);
                        
                        \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).this.parameter.Out.0\ <= \Quire Quire::op_Addition(Quire,UInt32).0.object2b25f3fa9b50e7492d78b34e15a583b8300db89f75b5c7cb2910bbab85a19ff0\;
                        \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).firstSegment.parameter.Out.0\ <= to_unsigned(1, 32);
                        \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).size.parameter.Out.0\ <= (\Quire Quire::op_Addition(Quire,UInt32).0.binaryOperationResult.0\);
                        \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Started.0\ <= true;
                        \Quire Quire::op_Addition(Quire,UInt32).0._State\ := \Quire Quire::op_Addition(Quire,UInt32).0._State_3\;
                        
                    when \Quire Quire::op_Addition(Quire,UInt32).0._State_3\ => 
                        
                        if (\Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Started.0\ = \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Finished.0\) then 
                            \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Started.0\ <= false;
                            \Quire Quire::op_Addition(Quire,UInt32).0.object2b25f3fa9b50e7492d78b34e15a583b8300db89f75b5c7cb2910bbab85a19ff0\ := \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).this.parameter.In.0\;
                            
                            
                            
                            
                            \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.Out.0\ <= \Quire Quire::op_Addition(Quire,UInt32).0.left\;
                            \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.Out.0\ <= \Quire Quire::op_Addition(Quire,UInt32).0.object2b25f3fa9b50e7492d78b34e15a583b8300db89f75b5c7cb2910bbab85a19ff0\;
                            \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\ <= true;
                            \Quire Quire::op_Addition(Quire,UInt32).0._State\ := \Quire Quire::op_Addition(Quire,UInt32).0._State_4\;
                        end if;
                        
                    when \Quire Quire::op_Addition(Quire,UInt32).0._State_4\ => 
                        
                        if (\Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\ = \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\) then 
                            \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\ <= false;
                            \Quire Quire::op_Addition(Quire,UInt32).0.return.0\ := \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).return.0\;
                            \Quire Quire::op_Addition(Quire,UInt32).0.left\ := \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.In.0\;
                            \Quire Quire::op_Addition(Quire,UInt32).0.object2b25f3fa9b50e7492d78b34e15a583b8300db89f75b5c7cb2910bbab85a19ff0\ := \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.In.0\;
                            \Quire Quire::op_Addition(Quire,UInt32).0.return\ <= \Quire Quire::op_Addition(Quire,UInt32).0.return.0\;
                            \Quire Quire::op_Addition(Quire,UInt32).0._State\ := \Quire Quire::op_Addition(Quire,UInt32).0._State_1\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Quire Quire::op_OnesComplement(Quire).0._StateMachine\: process (\Clock\) 
        Variable \Quire Quire::op_OnesComplement(Quire).0._State\: \Quire Quire::op_OnesComplement(Quire).0._States\ := \Quire Quire::op_OnesComplement(Quire).0._State_0\;
        Variable \Quire Quire::op_OnesComplement(Quire).0.q\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire Quire::op_OnesComplement(Quire).0.num\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_OnesComplement(Quire).0.binaryOperationResult.0\: boolean := false;
        Variable \Quire Quire::op_OnesComplement(Quire).0.unaryOperationResult.0\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_OnesComplement(Quire).0.binaryOperationResult.1\: unsigned(15 downto 0) := to_unsigned(0, 16);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Quire Quire::op_OnesComplement(Quire).0._Finished\ <= false;
                \Quire Quire::op_OnesComplement(Quire).0._State\ := \Quire Quire::op_OnesComplement(Quire).0._State_0\;
                \Quire Quire::op_OnesComplement(Quire).0.num\ := to_unsigned(0, 16);
                \Quire Quire::op_OnesComplement(Quire).0.binaryOperationResult.0\ := false;
                \Quire Quire::op_OnesComplement(Quire).0.unaryOperationResult.0\ := to_unsigned(0, 64);
                \Quire Quire::op_OnesComplement(Quire).0.binaryOperationResult.1\ := to_unsigned(0, 16);
            else 
                case \Quire Quire::op_OnesComplement(Quire).0._State\ is 
                    when \Quire Quire::op_OnesComplement(Quire).0._State_0\ => 
                        
                        
                        if (\Quire Quire::op_OnesComplement(Quire).0._Started\ = true) then 
                            \Quire Quire::op_OnesComplement(Quire).0._State\ := \Quire Quire::op_OnesComplement(Quire).0._State_2\;
                        end if;
                        
                    when \Quire Quire::op_OnesComplement(Quire).0._State_1\ => 
                        
                        
                        if (\Quire Quire::op_OnesComplement(Quire).0._Started\ = true) then 
                            \Quire Quire::op_OnesComplement(Quire).0._Finished\ <= true;
                        else 
                            \Quire Quire::op_OnesComplement(Quire).0._Finished\ <= false;
                            \Quire Quire::op_OnesComplement(Quire).0._State\ := \Quire Quire::op_OnesComplement(Quire).0._State_0\;
                        end if;
                        
                        \Quire Quire::op_OnesComplement(Quire).0.q.parameter.Out\ <= \Quire Quire::op_OnesComplement(Quire).0.q\;
                        
                    when \Quire Quire::op_OnesComplement(Quire).0._State_2\ => 
                        \Quire Quire::op_OnesComplement(Quire).0.q\ := \Quire Quire::op_OnesComplement(Quire).0.q.parameter.In\;
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_OnesComplement(Quire).0.num\ := SmartResize(unsigned(to_signed(0, 32)), 16);
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_OnesComplement(Quire).0._State\ := \Quire Quire::op_OnesComplement(Quire).0._State_3\;
                        
                    when \Quire Quire::op_OnesComplement(Quire).0._State_3\ => 
                        
                        
                        \Quire Quire::op_OnesComplement(Quire).0.binaryOperationResult.0\ := signed(SmartResize((\Quire Quire::op_OnesComplement(Quire).0.num\), 32)) < signed(SmartResize((\Quire Quire::op_OnesComplement(Quire).0.q\.\SegmentCount\), 32));
                        if (\Quire Quire::op_OnesComplement(Quire).0.binaryOperationResult.0\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Quire::op_OnesComplement(Quire).0.unaryOperationResult.0\ := not(\Quire Quire::op_OnesComplement(Quire).0.q\.\Segments\(to_integer(\Quire Quire::op_OnesComplement(Quire).0.num\)));
                            \Quire Quire::op_OnesComplement(Quire).0.q\.\Segments\(to_integer(\Quire Quire::op_OnesComplement(Quire).0.num\)) := \Quire Quire::op_OnesComplement(Quire).0.unaryOperationResult.0\;
                            
                            
                            
                            \Quire Quire::op_OnesComplement(Quire).0._State\ := \Quire Quire::op_OnesComplement(Quire).0._State_5\;
                        else 
                            \Quire Quire::op_OnesComplement(Quire).0._State\ := \Quire Quire::op_OnesComplement(Quire).0._State_4\;
                        end if;
                        
                    when \Quire Quire::op_OnesComplement(Quire).0._State_4\ => 
                        
                        
                        
                        
                        \Quire Quire::op_OnesComplement(Quire).0.return\ <= \Quire Quire::op_OnesComplement(Quire).0.q\;
                        \Quire Quire::op_OnesComplement(Quire).0._State\ := \Quire Quire::op_OnesComplement(Quire).0._State_1\;
                        
                    when \Quire Quire::op_OnesComplement(Quire).0._State_5\ => 
                        
                        \Quire Quire::op_OnesComplement(Quire).0.binaryOperationResult.1\ := SmartResize(unsigned(signed(SmartResize((\Quire Quire::op_OnesComplement(Quire).0.num\), 32)) + to_signed(1, 32)), 16);
                        \Quire Quire::op_OnesComplement(Quire).0.num\ := (\Quire Quire::op_OnesComplement(Quire).0.binaryOperationResult.1\);
                        
                        if (\Quire Quire::op_OnesComplement(Quire).0._State\ = \Quire Quire::op_OnesComplement(Quire).0._State_5\) then 
                            \Quire Quire::op_OnesComplement(Quire).0._State\ := \Quire Quire::op_OnesComplement(Quire).0._State_3\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Boolean Quire::op_Equality(Quire,Quire).0._StateMachine\: process (\Clock\) 
        Variable \Boolean Quire::op_Equality(Quire,Quire).0._State\: \Boolean Quire::op_Equality(Quire,Quire).0._States\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_0\;
        Variable \Boolean Quire::op_Equality(Quire,Quire).0.left\: \Lombiq.Arithmetics.Quire\;
        Variable \Boolean Quire::op_Equality(Quire,Quire).0.right\: \Lombiq.Arithmetics.Quire\;
        Variable \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.0\: boolean := false;
        Variable \Boolean Quire::op_Equality(Quire,Quire).0.num\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.1\: boolean := false;
        Variable \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.2\: boolean := false;
        Variable \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.3\: unsigned(15 downto 0) := to_unsigned(0, 16);
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Boolean Quire::op_Equality(Quire,Quire).0._Finished\ <= false;
                \Boolean Quire::op_Equality(Quire,Quire).0.return\ <= false;
                \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_0\;
                \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.0\ := false;
                \Boolean Quire::op_Equality(Quire,Quire).0.num\ := to_unsigned(0, 16);
                \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.1\ := false;
                \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.2\ := false;
                \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.3\ := to_unsigned(0, 16);
            else 
                case \Boolean Quire::op_Equality(Quire,Quire).0._State\ is 
                    when \Boolean Quire::op_Equality(Quire,Quire).0._State_0\ => 
                        
                        
                        if (\Boolean Quire::op_Equality(Quire,Quire).0._Started\ = true) then 
                            \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_2\;
                        end if;
                        
                    when \Boolean Quire::op_Equality(Quire,Quire).0._State_1\ => 
                        
                        
                        if (\Boolean Quire::op_Equality(Quire,Quire).0._Started\ = true) then 
                            \Boolean Quire::op_Equality(Quire,Quire).0._Finished\ <= true;
                        else 
                            \Boolean Quire::op_Equality(Quire,Quire).0._Finished\ <= false;
                            \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_0\;
                        end if;
                        
                        \Boolean Quire::op_Equality(Quire,Quire).0.left.parameter.Out\ <= \Boolean Quire::op_Equality(Quire,Quire).0.left\;
                        \Boolean Quire::op_Equality(Quire,Quire).0.right.parameter.Out\ <= \Boolean Quire::op_Equality(Quire,Quire).0.right\;
                        
                    when \Boolean Quire::op_Equality(Quire,Quire).0._State_2\ => 
                        \Boolean Quire::op_Equality(Quire,Quire).0.left\ := \Boolean Quire::op_Equality(Quire,Quire).0.left.parameter.In\;
                        \Boolean Quire::op_Equality(Quire,Quire).0.right\ := \Boolean Quire::op_Equality(Quire,Quire).0.right.parameter.In\;
                        
                        
                        
                        
                        
                        \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.0\ := signed(SmartResize((\Boolean Quire::op_Equality(Quire,Quire).0.left\.\SegmentCount\), 32)) /= signed(SmartResize((\Boolean Quire::op_Equality(Quire,Quire).0.right\.\SegmentCount\), 32));

                        
                        
                        

                        if (\Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.0\) then 
                            \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_4\;
                        else 
                            
                            \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_3\;
                        end if;
                        
                    when \Boolean Quire::op_Equality(Quire,Quire).0._State_3\ => 
                        
                        
                        
                        
                        
                        
                        
                        \Boolean Quire::op_Equality(Quire,Quire).0.num\ := SmartResize(unsigned(to_signed(0, 32)), 16);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_5\;
                        
                    when \Boolean Quire::op_Equality(Quire,Quire).0._State_4\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Boolean Quire::op_Equality(Quire,Quire).0.return\ <= false;
                        \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_1\;
                        
                        if (\Boolean Quire::op_Equality(Quire,Quire).0._State\ = \Boolean Quire::op_Equality(Quire,Quire).0._State_4\) then 
                            \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_3\;
                        end if;
                        
                    when \Boolean Quire::op_Equality(Quire,Quire).0._State_5\ => 
                        
                        
                        \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.1\ := signed(SmartResize((\Boolean Quire::op_Equality(Quire,Quire).0.num\), 32)) < signed(SmartResize((\Boolean Quire::op_Equality(Quire,Quire).0.left\.\SegmentCount\), 32));
                        if (\Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.1\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.2\ := \Boolean Quire::op_Equality(Quire,Quire).0.left\.\Segments\(to_integer(\Boolean Quire::op_Equality(Quire,Quire).0.num\)) /= \Boolean Quire::op_Equality(Quire,Quire).0.right\.\Segments\(to_integer(\Boolean Quire::op_Equality(Quire,Quire).0.num\));

                            
                            
                            

                            if (\Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.2\) then 
                                \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_8\;
                            else 
                                
                                \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_7\;
                            end if;
                        else 
                            \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_6\;
                        end if;
                        
                    when \Boolean Quire::op_Equality(Quire,Quire).0._State_6\ => 
                        
                        
                        
                        
                        \Boolean Quire::op_Equality(Quire,Quire).0.return\ <= true;
                        \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_1\;
                        
                    when \Boolean Quire::op_Equality(Quire,Quire).0._State_7\ => 
                        
                        
                        
                        
                        \Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.3\ := SmartResize(unsigned(signed(SmartResize((\Boolean Quire::op_Equality(Quire,Quire).0.num\), 32)) + to_signed(1, 32)), 16);
                        \Boolean Quire::op_Equality(Quire,Quire).0.num\ := (\Boolean Quire::op_Equality(Quire,Quire).0.binaryOperationResult.3\);
                        
                        if (\Boolean Quire::op_Equality(Quire,Quire).0._State\ = \Boolean Quire::op_Equality(Quire,Quire).0._State_7\) then 
                            \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_5\;
                        end if;
                        
                    when \Boolean Quire::op_Equality(Quire,Quire).0._State_8\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Boolean Quire::op_Equality(Quire,Quire).0.return\ <= false;
                        \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_1\;
                        
                        if (\Boolean Quire::op_Equality(Quire,Quire).0._State\ = \Boolean Quire::op_Equality(Quire,Quire).0._State_8\) then 
                            \Boolean Quire::op_Equality(Quire,Quire).0._State\ := \Boolean Quire::op_Equality(Quire,Quire).0._State_7\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Quire Quire::op_RightShift(Quire,Int32).0._StateMachine\: process (\Clock\) 
        Variable \Quire Quire::op_RightShift(Quire,Int32).0._State\: \Quire Quire::op_RightShift(Quire,Int32).0._States\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_0\;
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.left\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.right\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.1\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.2\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.3\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.num\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.array\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.num2\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.4\: boolean := false;
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.flag\: boolean := false;
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.num3\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.5\: boolean := false;
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.num4\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.6\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.flag2\: boolean := false;
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.7\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.8\: boolean := false;
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.9\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.10\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.11\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.12\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_RightShift(Quire,Int32).0.object157c924d312931f99624f9990346efe22383342001d9935b6c35c3ad8da224b8\: \Lombiq.Arithmetics.Quire\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Quire Quire::op_RightShift(Quire,Int32).0._Finished\ <= false;
                \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 64));
                \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= false;
                \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_0\;
                \Quire Quire::op_RightShift(Quire,Int32).0.right\ := to_signed(0, 32);
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.0\ := to_signed(0, 32);
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.1\ := to_signed(0, 32);
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.2\ := to_signed(0, 32);
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.3\ := to_signed(0, 32);
                \Quire Quire::op_RightShift(Quire,Int32).0.num\ := to_unsigned(0, 64);
                \Quire Quire::op_RightShift(Quire,Int32).0.array\ := (others => to_unsigned(0, 64));
                \Quire Quire::op_RightShift(Quire,Int32).0.num2\ := to_unsigned(0, 16);
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.4\ := false;
                \Quire Quire::op_RightShift(Quire,Int32).0.flag\ := false;
                \Quire Quire::op_RightShift(Quire,Int32).0.num3\ := to_unsigned(0, 16);
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.5\ := false;
                \Quire Quire::op_RightShift(Quire,Int32).0.num4\ := to_unsigned(0, 16);
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.6\ := to_unsigned(0, 16);
                \Quire Quire::op_RightShift(Quire,Int32).0.flag2\ := false;
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.7\ := to_unsigned(0, 64);
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.8\ := false;
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.9\ := to_unsigned(0, 64);
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.10\ := to_unsigned(0, 64);
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.11\ := to_unsigned(0, 16);
                \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.12\ := to_unsigned(0, 16);
            else 
                case \Quire Quire::op_RightShift(Quire,Int32).0._State\ is 
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_0\ => 
                        
                        
                        if (\Quire Quire::op_RightShift(Quire,Int32).0._Started\ = true) then 
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_2\;
                        end if;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_1\ => 
                        
                        
                        if (\Quire Quire::op_RightShift(Quire,Int32).0._Started\ = true) then 
                            \Quire Quire::op_RightShift(Quire,Int32).0._Finished\ <= true;
                        else 
                            \Quire Quire::op_RightShift(Quire,Int32).0._Finished\ <= false;
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_0\;
                        end if;
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.left.parameter.Out\ <= \Quire Quire::op_RightShift(Quire,Int32).0.left\;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_2\ => 
                        \Quire Quire::op_RightShift(Quire,Int32).0.left\ := \Quire Quire::op_RightShift(Quire,Int32).0.left.parameter.In\;
                        \Quire Quire::op_RightShift(Quire,Int32).0.right\ := \Quire Quire::op_RightShift(Quire,Int32).0.right.parameter.In\;
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.0\ := SmartResize(signed(SmartResize((\Quire Quire::op_RightShift(Quire,Int32).0.left\.\SegmentCount\), 32)) * to_signed(6, 32), 32);
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.1\ := shift_left(to_signed(1, 32), to_integer(unsigned(SmartResize(\Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.0\, 5))));
                        \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_3\;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_3\ => 
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.2\ := (\Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.1\) - to_signed(1, 32);
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.3\ := \Quire Quire::op_RightShift(Quire,Int32).0.right\ and (\Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.2\);
                        \Quire Quire::op_RightShift(Quire,Int32).0.right\ := \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.3\;
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.num\ := "1000000000000000000000000000000000000000000000000000000000000000";
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.array\ := (others => to_unsigned(0, 64));
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.array\ := \Quire Quire::op_RightShift(Quire,Int32).0.left\.\Segments\(0 to 7);
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.num2\ := SmartResize(unsigned(to_signed(0, 32)), 16);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_4\;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_4\ => 
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.4\ := signed(SmartResize((\Quire Quire::op_RightShift(Quire,Int32).0.num2\), 32)) < (\Quire Quire::op_RightShift(Quire,Int32).0.right\);
                        if (\Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.4\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Quire::op_RightShift(Quire,Int32).0.flag\ := false;
                            
                            
                            
                            
                            
                            
                            \Quire Quire::op_RightShift(Quire,Int32).0.num3\ := SmartResize(unsigned(to_signed(1, 32)), 16);
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_6\;
                        else 
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_5\;
                        end if;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_5\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.object157c924d312931f99624f9990346efe22383342001d9935b6c35c3ad8da224b8\.\IsNull\ := false;
                        \Quire Quire::op_RightShift(Quire,Int32).0.object157c924d312931f99624f9990346efe22383342001d9935b6c35c3ad8da224b8\.\Size\ := to_unsigned(0, 16);
                        \Quire Quire::op_RightShift(Quire,Int32).0.object157c924d312931f99624f9990346efe22383342001d9935b6c35c3ad8da224b8\.\SegmentCount\ := to_unsigned(0, 16);
                        \Quire Quire::op_RightShift(Quire,Int32).0.object157c924d312931f99624f9990346efe22383342001d9935b6c35c3ad8da224b8\.\Segments\ := (others => to_unsigned(0, 64));
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\ <= \Quire Quire::op_RightShift(Quire,Int32).0.object157c924d312931f99624f9990346efe22383342001d9935b6c35c3ad8da224b8\;
                        \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\ <= \Quire Quire::op_RightShift(Quire,Int32).0.array\;
                        \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\ <= SmartResize(unsigned(to_signed(0, 32)), 16);
                        \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= true;
                        \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_12\;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_6\ => 
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.5\ := signed(SmartResize((\Quire Quire::op_RightShift(Quire,Int32).0.num3\), 32)) <= to_signed(8, 32);
                        if (\Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.5\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.6\ := SmartResize(unsigned(to_signed(8, 32) - signed(SmartResize((\Quire Quire::op_RightShift(Quire,Int32).0.num3\), 32))), 16);
                            \Quire Quire::op_RightShift(Quire,Int32).0.num4\ := (\Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.6\);
                            
                            
                            
                            
                            
                            
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_8\;
                        else 
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_7\;
                        end if;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_7\ => 
                        
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.12\ := SmartResize(unsigned(signed(SmartResize((\Quire Quire::op_RightShift(Quire,Int32).0.num2\), 32)) + to_signed(1, 32)), 16);
                        \Quire Quire::op_RightShift(Quire,Int32).0.num2\ := (\Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.12\);
                        
                        if (\Quire Quire::op_RightShift(Quire,Int32).0._State\ = \Quire Quire::op_RightShift(Quire,Int32).0._State_7\) then 
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_4\;
                        end if;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_8\ => 
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.7\ := \Quire Quire::op_RightShift(Quire,Int32).0.array\(to_integer(\Quire Quire::op_RightShift(Quire,Int32).0.num4\)) and to_unsigned(1, 64);
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.8\ := (\Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.7\) = to_unsigned(1, 64);
                        \Quire Quire::op_RightShift(Quire,Int32).0.flag2\ := \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.8\;
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_9\;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_9\ => 
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.9\ := SmartResize(shift_right(\Quire Quire::op_RightShift(Quire,Int32).0.array\(to_integer(\Quire Quire::op_RightShift(Quire,Int32).0.num4\)), to_integer(unsigned(SmartResize(to_signed(1, 32), 6) and "111111"))), 64);
                        \Quire Quire::op_RightShift(Quire,Int32).0.array\(to_integer(\Quire Quire::op_RightShift(Quire,Int32).0.num4\)) := \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.9\;
                        
                        
                        
                        
                        

                        
                        
                        

                        if (\Quire Quire::op_RightShift(Quire,Int32).0.flag\) then 
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_11\;
                        else 
                            
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_10\;
                        end if;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_10\ => 
                        
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.flag\ := \Quire Quire::op_RightShift(Quire,Int32).0.flag2\;
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.11\ := SmartResize(unsigned(signed(SmartResize((\Quire Quire::op_RightShift(Quire,Int32).0.num3\), 32)) + to_signed(1, 32)), 16);
                        \Quire Quire::op_RightShift(Quire,Int32).0.num3\ := (\Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.11\);
                        
                        if (\Quire Quire::op_RightShift(Quire,Int32).0._State\ = \Quire Quire::op_RightShift(Quire,Int32).0._State_10\) then 
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_6\;
                        end if;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_11\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.10\ := \Quire Quire::op_RightShift(Quire,Int32).0.array\(to_integer(\Quire Quire::op_RightShift(Quire,Int32).0.num4\)) or \Quire Quire::op_RightShift(Quire,Int32).0.num\;
                        \Quire Quire::op_RightShift(Quire,Int32).0.array\(to_integer(\Quire Quire::op_RightShift(Quire,Int32).0.num4\)) := \Quire Quire::op_RightShift(Quire,Int32).0.binaryOperationResult.10\;
                        
                        if (\Quire Quire::op_RightShift(Quire,Int32).0._State\ = \Quire Quire::op_RightShift(Quire,Int32).0._State_11\) then 
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_10\;
                        end if;
                        
                    when \Quire Quire::op_RightShift(Quire,Int32).0._State_12\ => 
                        
                        if (\Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ = \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\) then 
                            \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= false;
                            \Quire Quire::op_RightShift(Quire,Int32).0.object157c924d312931f99624f9990346efe22383342001d9935b6c35c3ad8da224b8\ := \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\;
                            \Quire Quire::op_RightShift(Quire,Int32).0.array\ := \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\;
                            
                            
                            
                            \Quire Quire::op_RightShift(Quire,Int32).0.return\ <= \Quire Quire::op_RightShift(Quire,Int32).0.object157c924d312931f99624f9990346efe22383342001d9935b6c35c3ad8da224b8\;
                            \Quire Quire::op_RightShift(Quire,Int32).0._State\ := \Quire Quire::op_RightShift(Quire,Int32).0._State_1\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Quire Quire::op_LeftShift(Quire,Int32).0._StateMachine\: process (\Clock\) 
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0._State\: \Quire Quire::op_LeftShift(Quire,Int32).0._States\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_0\;
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.left\: \Lombiq.Arithmetics.Quire\;
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.right\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.0\: signed(31 downto 0) := to_signed(0, 32);
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.num\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.array\: \unsigned64_Array\(0 to 7) := (others => to_unsigned(0, 64));
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.num2\: unsigned(31 downto 0) := to_unsigned(0, 32);
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.num3\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.1\: boolean := false;
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.flag\: boolean := false;
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.num4\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.2\: boolean := false;
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.flag2\: boolean := false;
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.3\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.4\: boolean := false;
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.5\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.6\: unsigned(63 downto 0) := to_unsigned(0, 64);
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.7\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.8\: unsigned(15 downto 0) := to_unsigned(0, 16);
        Variable \Quire Quire::op_LeftShift(Quire,Int32).0.objectc996901721b3380940539d5e2ccc153d36bc5159fbc7657e5cc431d1b5e93c1f\: \Lombiq.Arithmetics.Quire\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Quire Quire::op_LeftShift(Quire,Int32).0._Finished\ <= false;
                \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\ <= (others => to_unsigned(0, 64));
                \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\ <= to_unsigned(0, 16);
                \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= false;
                \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_0\;
                \Quire Quire::op_LeftShift(Quire,Int32).0.right\ := to_signed(0, 32);
                \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.0\ := to_signed(0, 32);
                \Quire Quire::op_LeftShift(Quire,Int32).0.num\ := to_unsigned(0, 64);
                \Quire Quire::op_LeftShift(Quire,Int32).0.array\ := (others => to_unsigned(0, 64));
                \Quire Quire::op_LeftShift(Quire,Int32).0.num2\ := to_unsigned(0, 32);
                \Quire Quire::op_LeftShift(Quire,Int32).0.num3\ := to_unsigned(0, 16);
                \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.1\ := false;
                \Quire Quire::op_LeftShift(Quire,Int32).0.flag\ := false;
                \Quire Quire::op_LeftShift(Quire,Int32).0.num4\ := to_unsigned(0, 16);
                \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.2\ := false;
                \Quire Quire::op_LeftShift(Quire,Int32).0.flag2\ := false;
                \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.3\ := to_unsigned(0, 64);
                \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.4\ := false;
                \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.5\ := to_unsigned(0, 64);
                \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.6\ := to_unsigned(0, 64);
                \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.7\ := to_unsigned(0, 16);
                \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.8\ := to_unsigned(0, 16);
            else 
                case \Quire Quire::op_LeftShift(Quire,Int32).0._State\ is 
                    when \Quire Quire::op_LeftShift(Quire,Int32).0._State_0\ => 
                        
                        
                        if (\Quire Quire::op_LeftShift(Quire,Int32).0._Started\ = true) then 
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_2\;
                        end if;
                        
                    when \Quire Quire::op_LeftShift(Quire,Int32).0._State_1\ => 
                        
                        
                        if (\Quire Quire::op_LeftShift(Quire,Int32).0._Started\ = true) then 
                            \Quire Quire::op_LeftShift(Quire,Int32).0._Finished\ <= true;
                        else 
                            \Quire Quire::op_LeftShift(Quire,Int32).0._Finished\ <= false;
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_0\;
                        end if;
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.left.parameter.Out\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.left\;
                        
                    when \Quire Quire::op_LeftShift(Quire,Int32).0._State_2\ => 
                        \Quire Quire::op_LeftShift(Quire,Int32).0.left\ := \Quire Quire::op_LeftShift(Quire,Int32).0.left.parameter.In\;
                        \Quire Quire::op_LeftShift(Quire,Int32).0.right\ := \Quire Quire::op_LeftShift(Quire,Int32).0.right.parameter.In\;
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.0\ := \Quire Quire::op_LeftShift(Quire,Int32).0.right\ and to_signed(65535, 32);
                        \Quire Quire::op_LeftShift(Quire,Int32).0.right\ := \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.0\;
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.num\ := "1000000000000000000000000000000000000000000000000000000000000000";
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.array\ := (others => to_unsigned(0, 64));
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.array\ := \Quire Quire::op_LeftShift(Quire,Int32).0.left\.\Segments\(0 to 7);
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.num2\ := to_unsigned(1, 32);
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.num3\ := SmartResize(unsigned(to_signed(0, 32)), 16);
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_3\;
                        
                    when \Quire Quire::op_LeftShift(Quire,Int32).0._State_3\ => 
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.1\ := signed(SmartResize((\Quire Quire::op_LeftShift(Quire,Int32).0.num3\), 32)) < (\Quire Quire::op_LeftShift(Quire,Int32).0.right\);
                        if (\Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.1\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Quire::op_LeftShift(Quire,Int32).0.flag\ := false;
                            
                            
                            
                            
                            
                            
                            \Quire Quire::op_LeftShift(Quire,Int32).0.num4\ := SmartResize(unsigned(to_signed(0, 32)), 16);
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_5\;
                        else 
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_4\;
                        end if;
                        
                    when \Quire Quire::op_LeftShift(Quire,Int32).0._State_4\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.objectc996901721b3380940539d5e2ccc153d36bc5159fbc7657e5cc431d1b5e93c1f\.\IsNull\ := false;
                        \Quire Quire::op_LeftShift(Quire,Int32).0.objectc996901721b3380940539d5e2ccc153d36bc5159fbc7657e5cc431d1b5e93c1f\.\Size\ := to_unsigned(0, 16);
                        \Quire Quire::op_LeftShift(Quire,Int32).0.objectc996901721b3380940539d5e2ccc153d36bc5159fbc7657e5cc431d1b5e93c1f\.\SegmentCount\ := to_unsigned(0, 16);
                        \Quire Quire::op_LeftShift(Quire,Int32).0.objectc996901721b3380940539d5e2ccc153d36bc5159fbc7657e5cc431d1b5e93c1f\.\Segments\ := (others => to_unsigned(0, 64));
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.objectc996901721b3380940539d5e2ccc153d36bc5159fbc7657e5cc431d1b5e93c1f\;
                        \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.array\;
                        \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\ <= SmartResize(unsigned(to_signed(0, 32)), 16);
                        \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= true;
                        \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_10\;
                        
                    when \Quire Quire::op_LeftShift(Quire,Int32).0._State_5\ => 
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.2\ := signed(SmartResize((\Quire Quire::op_LeftShift(Quire,Int32).0.num4\), 32)) < to_signed(8, 32);
                        if (\Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.2\) then 
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            
                            \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.3\ := \Quire Quire::op_LeftShift(Quire,Int32).0.array\(to_integer(\Quire Quire::op_LeftShift(Quire,Int32).0.num4\)) and \Quire Quire::op_LeftShift(Quire,Int32).0.num\;
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_7\;
                        else 
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_6\;
                        end if;
                        
                    when \Quire Quire::op_LeftShift(Quire,Int32).0._State_6\ => 
                        
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.8\ := SmartResize(unsigned(signed(SmartResize((\Quire Quire::op_LeftShift(Quire,Int32).0.num3\), 32)) + to_signed(1, 32)), 16);
                        \Quire Quire::op_LeftShift(Quire,Int32).0.num3\ := (\Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.8\);
                        
                        if (\Quire Quire::op_LeftShift(Quire,Int32).0._State\ = \Quire Quire::op_LeftShift(Quire,Int32).0._State_6\) then 
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_3\;
                        end if;
                        
                    when \Quire Quire::op_LeftShift(Quire,Int32).0._State_7\ => 
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.4\ := (\Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.3\) = \Quire Quire::op_LeftShift(Quire,Int32).0.num\;
                        \Quire Quire::op_LeftShift(Quire,Int32).0.flag2\ := \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.4\;
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.5\ := SmartResize(shift_left(\Quire Quire::op_LeftShift(Quire,Int32).0.array\(to_integer(\Quire Quire::op_LeftShift(Quire,Int32).0.num4\)), to_integer(unsigned(SmartResize(to_signed(1, 32), 6)))), 64);
                        \Quire Quire::op_LeftShift(Quire,Int32).0.array\(to_integer(\Quire Quire::op_LeftShift(Quire,Int32).0.num4\)) := \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.5\;
                        
                        
                        
                        
                        

                        
                        
                        

                        if (\Quire Quire::op_LeftShift(Quire,Int32).0.flag\) then 
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_9\;
                        else 
                            
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_8\;
                        end if;
                        
                    when \Quire Quire::op_LeftShift(Quire,Int32).0._State_8\ => 
                        
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.flag\ := \Quire Quire::op_LeftShift(Quire,Int32).0.flag2\;
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.7\ := SmartResize(unsigned(signed(SmartResize((\Quire Quire::op_LeftShift(Quire,Int32).0.num4\), 32)) + to_signed(1, 32)), 16);
                        \Quire Quire::op_LeftShift(Quire,Int32).0.num4\ := (\Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.7\);
                        
                        if (\Quire Quire::op_LeftShift(Quire,Int32).0._State\ = \Quire Quire::op_LeftShift(Quire,Int32).0._State_8\) then 
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_5\;
                        end if;
                        
                    when \Quire Quire::op_LeftShift(Quire,Int32).0._State_9\ => 
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        \Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.6\ := \Quire Quire::op_LeftShift(Quire,Int32).0.array\(to_integer(\Quire Quire::op_LeftShift(Quire,Int32).0.num4\)) or SmartResize((\Quire Quire::op_LeftShift(Quire,Int32).0.num2\), 64);
                        \Quire Quire::op_LeftShift(Quire,Int32).0.array\(to_integer(\Quire Quire::op_LeftShift(Quire,Int32).0.num4\)) := (\Quire Quire::op_LeftShift(Quire,Int32).0.binaryOperationResult.6\);
                        
                        if (\Quire Quire::op_LeftShift(Quire,Int32).0._State\ = \Quire Quire::op_LeftShift(Quire,Int32).0._State_9\) then 
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_8\;
                        end if;
                        
                    when \Quire Quire::op_LeftShift(Quire,Int32).0._State_10\ => 
                        
                        if (\Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ = \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\) then 
                            \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ <= false;
                            \Quire Quire::op_LeftShift(Quire,Int32).0.objectc996901721b3380940539d5e2ccc153d36bc5159fbc7657e5cc431d1b5e93c1f\ := \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\;
                            \Quire Quire::op_LeftShift(Quire,Int32).0.array\ := \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\;
                            
                            
                            
                            \Quire Quire::op_LeftShift(Quire,Int32).0.return\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.objectc996901721b3380940539d5e2ccc153d36bc5159fbc7657e5cc431d1b5e93c1f\;
                            \Quire Quire::op_LeftShift(Quire,Int32).0._State\ := \Quire Quire::op_LeftShift(Quire,Int32).0._State_1\;
                        end if;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \UInt64 Quire::op_Explicit(Quire).0._StateMachine\: process (\Clock\) 
        Variable \UInt64 Quire::op_Explicit(Quire).0._State\: \UInt64 Quire::op_Explicit(Quire).0._States\ := \UInt64 Quire::op_Explicit(Quire).0._State_0\;
        Variable \UInt64 Quire::op_Explicit(Quire).0.x\: \Lombiq.Arithmetics.Quire\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \UInt64 Quire::op_Explicit(Quire).0._Finished\ <= false;
                \UInt64 Quire::op_Explicit(Quire).0.return\ <= to_unsigned(0, 64);
                \UInt64 Quire::op_Explicit(Quire).0._State\ := \UInt64 Quire::op_Explicit(Quire).0._State_0\;
            else 
                case \UInt64 Quire::op_Explicit(Quire).0._State\ is 
                    when \UInt64 Quire::op_Explicit(Quire).0._State_0\ => 
                        
                        
                        if (\UInt64 Quire::op_Explicit(Quire).0._Started\ = true) then 
                            \UInt64 Quire::op_Explicit(Quire).0._State\ := \UInt64 Quire::op_Explicit(Quire).0._State_2\;
                        end if;
                        
                    when \UInt64 Quire::op_Explicit(Quire).0._State_1\ => 
                        
                        
                        if (\UInt64 Quire::op_Explicit(Quire).0._Started\ = true) then 
                            \UInt64 Quire::op_Explicit(Quire).0._Finished\ <= true;
                        else 
                            \UInt64 Quire::op_Explicit(Quire).0._Finished\ <= false;
                            \UInt64 Quire::op_Explicit(Quire).0._State\ := \UInt64 Quire::op_Explicit(Quire).0._State_0\;
                        end if;
                        
                        \UInt64 Quire::op_Explicit(Quire).0.x.parameter.Out\ <= \UInt64 Quire::op_Explicit(Quire).0.x\;
                        
                    when \UInt64 Quire::op_Explicit(Quire).0._State_2\ => 
                        \UInt64 Quire::op_Explicit(Quire).0.x\ := \UInt64 Quire::op_Explicit(Quire).0.x.parameter.In\;
                        
                        
                        
                        \UInt64 Quire::op_Explicit(Quire).0.return\ <= \UInt64 Quire::op_Explicit(Quire).0.x\.\Segments\(to_integer(to_signed(0, 32)));
                        \UInt64 Quire::op_Explicit(Quire).0._State\ := \UInt64 Quire::op_Explicit(Quire).0._State_1\;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \UInt32 Quire::op_Explicit(Quire).0._StateMachine\: process (\Clock\) 
        Variable \UInt32 Quire::op_Explicit(Quire).0._State\: \UInt32 Quire::op_Explicit(Quire).0._States\ := \UInt32 Quire::op_Explicit(Quire).0._State_0\;
        Variable \UInt32 Quire::op_Explicit(Quire).0.x\: \Lombiq.Arithmetics.Quire\;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \UInt32 Quire::op_Explicit(Quire).0._Finished\ <= false;
                \UInt32 Quire::op_Explicit(Quire).0.return\ <= to_unsigned(0, 32);
                \UInt32 Quire::op_Explicit(Quire).0._State\ := \UInt32 Quire::op_Explicit(Quire).0._State_0\;
            else 
                case \UInt32 Quire::op_Explicit(Quire).0._State\ is 
                    when \UInt32 Quire::op_Explicit(Quire).0._State_0\ => 
                        
                        
                        if (\UInt32 Quire::op_Explicit(Quire).0._Started\ = true) then 
                            \UInt32 Quire::op_Explicit(Quire).0._State\ := \UInt32 Quire::op_Explicit(Quire).0._State_2\;
                        end if;
                        
                    when \UInt32 Quire::op_Explicit(Quire).0._State_1\ => 
                        
                        
                        if (\UInt32 Quire::op_Explicit(Quire).0._Started\ = true) then 
                            \UInt32 Quire::op_Explicit(Quire).0._Finished\ <= true;
                        else 
                            \UInt32 Quire::op_Explicit(Quire).0._Finished\ <= false;
                            \UInt32 Quire::op_Explicit(Quire).0._State\ := \UInt32 Quire::op_Explicit(Quire).0._State_0\;
                        end if;
                        
                        \UInt32 Quire::op_Explicit(Quire).0.x.parameter.Out\ <= \UInt32 Quire::op_Explicit(Quire).0.x\;
                        
                    when \UInt32 Quire::op_Explicit(Quire).0._State_2\ => 
                        \UInt32 Quire::op_Explicit(Quire).0.x\ := \UInt32 Quire::op_Explicit(Quire).0.x.parameter.In\;
                        
                        
                        
                        \UInt32 Quire::op_Explicit(Quire).0.return\ <= SmartResize(\UInt32 Quire::op_Explicit(Quire).0.x\.\Segments\(to_integer(to_signed(0, 32))), 32);
                        \UInt32 Quire::op_Explicit(Quire).0._State\ := \UInt32 Quire::op_Explicit(Quire).0._State_1\;
                        
                end case;
            end if;
        end if;
    end process;
    


    
    \Finished\ <= \FinishedInternal\;
    \Hast::ExternalInvocationProxy()\: process (\Clock\) 
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \FinishedInternal\ <= false;
                \Hast::ExternalInvocationProxy().Posit32FusedCalculator::CalculateFusedSum(SimpleMemory)._Started.0\ <= false;
            else 
                if (\Started\ = true and \FinishedInternal\ = false) then 
                    
                    case \MemberId\ is 
                        when 0 => 
                            if (\Hast::ExternalInvocationProxy().Posit32FusedCalculator::CalculateFusedSum(SimpleMemory)._Started.0\ = false) then 
                                \Hast::ExternalInvocationProxy().Posit32FusedCalculator::CalculateFusedSum(SimpleMemory)._Started.0\ <= true;
                            elsif (\Hast::ExternalInvocationProxy().Posit32FusedCalculator::CalculateFusedSum(SimpleMemory)._Started.0\ = \Hast::ExternalInvocationProxy().Posit32FusedCalculator::CalculateFusedSum(SimpleMemory)._Finished.0\) then 
                                \Hast::ExternalInvocationProxy().Posit32FusedCalculator::CalculateFusedSum(SimpleMemory)._Started.0\ <= false;
                                \FinishedInternal\ <= true;
                            end if;
                        when others => 
                            null;
                    end case;
                else 
                    
                    if (\Started\ = false and \FinishedInternal\ = true) then 
                        \FinishedInternal\ <= false;
                    end if;
                end if;
            end if;
        end if;
    end process;
    


    
    
    \Posit32::.ctor(Int32).0._Started\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Started.0\;
    \Posit32::.ctor(Int32).0.this.parameter.In\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).this.parameter.Out.0\;
    \Posit32::.ctor(Int32).0.value.parameter.In\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).value.parameter.Out.0\;
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32)._Finished.0\ <= \Posit32::.ctor(Int32).0._Finished\;
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Int32).this.parameter.In.0\ <= \Posit32::.ctor(Int32).0.this.parameter.Out\;
    


    
    \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForStarted;
                \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\ <= false;
                \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\ <= false;
            else 

                
                case \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Started.0\) then 
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.runningIndex.0\ := 0;
                            \Quire Posit32::op_Explicit(Posit32).0._Started\ <= true;
                            \Quire Posit32::op_Explicit(Posit32).0.x.parameter.In\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32).x.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire Posit32::op_Explicit(Posit32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.runningState.0\ := AfterFinished;
                                    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\ <= true;
                                    \Quire Posit32::op_Explicit(Posit32).0._Started\ <= false;
                                    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32).return.0\ <= \Quire Posit32::op_Explicit(Posit32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.runningState.0\ := WaitingForStarted;
                            \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Started.0\) then 
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ := 0;
                            \Quire Posit32::op_Explicit(Posit32).0._Started\ <= true;
                            \Quire Posit32::op_Explicit(Posit32).0.x.parameter.In\ <= \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32).x.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire Posit32::op_Explicit(Posit32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := AfterFinished;
                                    \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\ <= true;
                                    \Quire Posit32::op_Explicit(Posit32).0._Started\ <= false;
                                    \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32).return.0\ <= \Quire Posit32::op_Explicit(Posit32).0.return\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire Posit32::op_Explicit(Posit32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForStarted;
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Posit32::op_Explicit(Posit32)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    


    
    
    \Posit32::.ctor(UInt32,Boolean).0._Started\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean)._Started.0\;
    \Posit32::.ctor(UInt32,Boolean).0.this.parameter.In\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).this.parameter.Out.0\;
    \Posit32::.ctor(UInt32,Boolean).0.bits.parameter.In\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).bits.parameter.Out.0\;
    \Posit32::.ctor(UInt32,Boolean).0.fromBitMask.parameter.In\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).fromBitMask.parameter.Out.0\;
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean)._Finished.0\ <= \Posit32::.ctor(UInt32,Boolean).0._Finished\;
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(UInt32,Boolean).this.parameter.In.0\ <= \Posit32::.ctor(UInt32,Boolean).0.this.parameter.Out\;
    


    
    
    \Posit32::FusedSum(Posit32[],Quire).0._Started\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire)._Started.0\;
    \Posit32::FusedSum(Posit32[],Quire).0.posits.parameter.In\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).posits.parameter.Out.0\;
    \Posit32::FusedSum(Posit32[],Quire).0.startingValue.parameter.In\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).startingValue.parameter.Out.0\;
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire)._Finished.0\ <= \Posit32::FusedSum(Posit32[],Quire).0._Finished\;
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).return.0\ <= \Posit32::FusedSum(Posit32[],Quire).0.return\;
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).posits.parameter.In.0\ <= \Posit32::FusedSum(Posit32[],Quire).0.posits.parameter.Out\;
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::FusedSum(Posit32[],Quire).startingValue.parameter.In.0\ <= \Posit32::FusedSum(Posit32[],Quire).0.startingValue.parameter.Out\;
    


    
    
    \Posit32::.ctor(Quire).0._Started\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire)._Started.0\;
    \Posit32::.ctor(Quire).0.this.parameter.In\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).this.parameter.Out.0\;
    \Posit32::.ctor(Quire).0.q.parameter.In\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).q.parameter.Out.0\;
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire)._Finished.0\ <= \Posit32::.ctor(Quire).0._Finished\;
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).this.parameter.In.0\ <= \Posit32::.ctor(Quire).0.this.parameter.Out\;
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.Posit32::.ctor(Quire).q.parameter.In.0\ <= \Posit32::.ctor(Quire).0.q.parameter.Out\;
    


    
    
    \Quire Quire::op_RightShift(Quire,Int32).0._Started\ <= \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Started.0\;
    \Quire Quire::op_RightShift(Quire,Int32).0.left.parameter.In\ <= \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.Out.0\;
    \Quire Quire::op_RightShift(Quire,Int32).0.right.parameter.In\ <= \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).right.parameter.Out.0\;
    \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32)._Finished.0\ <= \Quire Quire::op_RightShift(Quire,Int32).0._Finished\;
    \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).return.0\ <= \Quire Quire::op_RightShift(Quire,Int32).0.return\;
    \Posit32::.ctor(Quire).0.Quire Quire::op_RightShift(Quire,Int32).left.parameter.In.0\ <= \Quire Quire::op_RightShift(Quire,Int32).0.left.parameter.Out\;
    


    
    
    \UInt64 Quire::op_Explicit(Quire).0._Started\ <= \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Started.0\;
    \UInt64 Quire::op_Explicit(Quire).0.x.parameter.In\ <= \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).x.parameter.Out.0\;
    \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire)._Finished.0\ <= \UInt64 Quire::op_Explicit(Quire).0._Finished\;
    \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).return.0\ <= \UInt64 Quire::op_Explicit(Quire).0.return\;
    \Posit32::.ctor(Quire).0.UInt64 Quire::op_Explicit(Quire).x.parameter.In.0\ <= \UInt64 Quire::op_Explicit(Quire).0.x.parameter.Out\;
    


    
    \Hast::InternalInvocationProxy().Quire Quire::op_OnesComplement(Quire)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_OnesComplement(Quire).Posit32::.ctor(Quire).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_OnesComplement(Quire).Posit32::.ctor(Quire).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_OnesComplement(Quire).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_OnesComplement(Quire).Quire Posit32::op_Explicit(Posit32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Hast::InternalInvocationProxy().Quire Quire::op_OnesComplement(Quire).Posit32::.ctor(Quire).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire Quire::op_OnesComplement(Quire).Posit32::.ctor(Quire).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Quire Quire::op_OnesComplement(Quire).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire Quire::op_OnesComplement(Quire).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForStarted;
                \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire)._Finished.0\ <= false;
                \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_OnesComplement(Quire)._Finished.0\ <= false;
            else 

                
                case \Hast::InternalInvocationProxy().Quire Quire::op_OnesComplement(Quire).Posit32::.ctor(Quire).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire)._Started.0\) then 
                            \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire Quire::op_OnesComplement(Quire).Posit32::.ctor(Quire).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire Quire::op_OnesComplement(Quire).Posit32::.ctor(Quire).0.runningIndex.0\ := 0;
                            \Quire Quire::op_OnesComplement(Quire).0._Started\ <= true;
                            \Quire Quire::op_OnesComplement(Quire).0.q.parameter.In\ <= \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire).q.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire Quire::op_OnesComplement(Quire).Posit32::.ctor(Quire).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire Quire::op_OnesComplement(Quire).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire Quire::op_OnesComplement(Quire).Posit32::.ctor(Quire).0.runningState.0\ := AfterFinished;
                                    \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire)._Finished.0\ <= true;
                                    \Quire Quire::op_OnesComplement(Quire).0._Started\ <= false;
                                    \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire).return.0\ <= \Quire Quire::op_OnesComplement(Quire).0.return\;
                                    \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire).q.parameter.In.0\ <= \Quire Quire::op_OnesComplement(Quire).0.q.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire Quire::op_OnesComplement(Quire).Posit32::.ctor(Quire).0.runningState.0\ := WaitingForStarted;
                            \Posit32::.ctor(Quire).0.Quire Quire::op_OnesComplement(Quire)._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Quire Quire::op_OnesComplement(Quire).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_OnesComplement(Quire)._Started.0\) then 
                            \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_OnesComplement(Quire)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire Quire::op_OnesComplement(Quire).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire Quire::op_OnesComplement(Quire).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ := 0;
                            \Quire Quire::op_OnesComplement(Quire).0._Started\ <= true;
                            \Quire Quire::op_OnesComplement(Quire).0.q.parameter.In\ <= \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_OnesComplement(Quire).q.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire Quire::op_OnesComplement(Quire).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire Quire::op_OnesComplement(Quire).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire Quire::op_OnesComplement(Quire).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := AfterFinished;
                                    \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_OnesComplement(Quire)._Finished.0\ <= true;
                                    \Quire Quire::op_OnesComplement(Quire).0._Started\ <= false;
                                    \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_OnesComplement(Quire).return.0\ <= \Quire Quire::op_OnesComplement(Quire).0.return\;
                                    \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_OnesComplement(Quire).q.parameter.In.0\ <= \Quire Quire::op_OnesComplement(Quire).0.q.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_OnesComplement(Quire)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire Quire::op_OnesComplement(Quire).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForStarted;
                            \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_OnesComplement(Quire)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    


    
    \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,UInt32)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,UInt32).Posit32::.ctor(Quire).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,UInt32).Posit32::.ctor(Quire).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,UInt32).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,UInt32).Quire Posit32::op_Explicit(Posit32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,UInt32).Posit32::.ctor(Quire).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,UInt32).Posit32::.ctor(Quire).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,UInt32).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,UInt32).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForStarted;
                \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32)._Finished.0\ <= false;
                \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32)._Finished.0\ <= false;
            else 

                
                case \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,UInt32).Posit32::.ctor(Quire).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32)._Started.0\) then 
                            \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,UInt32).Posit32::.ctor(Quire).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,UInt32).Posit32::.ctor(Quire).0.runningIndex.0\ := 0;
                            \Quire Quire::op_Addition(Quire,UInt32).0._Started\ <= true;
                            \Quire Quire::op_Addition(Quire,UInt32).0.left.parameter.In\ <= \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).left.parameter.Out.0\;
                            \Quire Quire::op_Addition(Quire,UInt32).0.right.parameter.In\ <= \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,UInt32).Posit32::.ctor(Quire).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire Quire::op_Addition(Quire,UInt32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,UInt32).Posit32::.ctor(Quire).0.runningState.0\ := AfterFinished;
                                    \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32)._Finished.0\ <= true;
                                    \Quire Quire::op_Addition(Quire,UInt32).0._Started\ <= false;
                                    \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).return.0\ <= \Quire Quire::op_Addition(Quire,UInt32).0.return\;
                                    \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32).left.parameter.In.0\ <= \Quire Quire::op_Addition(Quire,UInt32).0.left.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,UInt32).Posit32::.ctor(Quire).0.runningState.0\ := WaitingForStarted;
                            \Posit32::.ctor(Quire).0.Quire Quire::op_Addition(Quire,UInt32)._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,UInt32).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32)._Started.0\) then 
                            \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,UInt32).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,UInt32).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ := 0;
                            \Quire Quire::op_Addition(Quire,UInt32).0._Started\ <= true;
                            \Quire Quire::op_Addition(Quire,UInt32).0.left.parameter.In\ <= \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32).left.parameter.Out.0\;
                            \Quire Quire::op_Addition(Quire,UInt32).0.right.parameter.In\ <= \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,UInt32).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire Quire::op_Addition(Quire,UInt32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,UInt32).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := AfterFinished;
                                    \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32)._Finished.0\ <= true;
                                    \Quire Quire::op_Addition(Quire,UInt32).0._Started\ <= false;
                                    \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32).return.0\ <= \Quire Quire::op_Addition(Quire,UInt32).0.return\;
                                    \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32).left.parameter.In.0\ <= \Quire Quire::op_Addition(Quire,UInt32).0.left.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,UInt32).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForStarted;
                            \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_Addition(Quire,UInt32)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    


    
    \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::.ctor(Quire).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::.ctor(Quire).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Quire Posit32::op_Explicit(Posit32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::.ctor(Quire).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::.ctor(Quire).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForStarted;
                \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= false;
                \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= false;
                \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= false;
            else 

                
                case \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::.ctor(Quire).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\) then 
                            \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::.ctor(Quire).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::.ctor(Quire).0.runningIndex.0\ := 0;
                            \Quire Quire::op_LeftShift(Quire,Int32).0._Started\ <= true;
                            \Quire Quire::op_LeftShift(Quire,Int32).0.left.parameter.In\ <= \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.Out.0\;
                            \Quire Quire::op_LeftShift(Quire,Int32).0.right.parameter.In\ <= \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::.ctor(Quire).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire Quire::op_LeftShift(Quire,Int32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::.ctor(Quire).0.runningState.0\ := AfterFinished;
                                    \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= true;
                                    \Quire Quire::op_LeftShift(Quire,Int32).0._Started\ <= false;
                                    \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).return.0\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.return\;
                                    \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.In.0\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.left.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::.ctor(Quire).0.runningState.0\ := WaitingForStarted;
                            \Posit32::.ctor(Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\) then 
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ := 0;
                            \Quire Quire::op_LeftShift(Quire,Int32).0._Started\ <= true;
                            \Quire Quire::op_LeftShift(Quire,Int32).0.left.parameter.In\ <= \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.Out.0\;
                            \Quire Quire::op_LeftShift(Quire,Int32).0.right.parameter.In\ <= \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire Quire::op_LeftShift(Quire,Int32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := AfterFinished;
                                    \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= true;
                                    \Quire Quire::op_LeftShift(Quire,Int32).0._Started\ <= false;
                                    \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).return.0\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.return\;
                                    \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.In.0\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.left.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForStarted;
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\) then 
                            \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ := 0;
                            \Quire Quire::op_LeftShift(Quire,Int32).0._Started\ <= true;
                            \Quire Quire::op_LeftShift(Quire,Int32).0.left.parameter.In\ <= \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.Out.0\;
                            \Quire Quire::op_LeftShift(Quire,Int32).0.right.parameter.In\ <= \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire Quire::op_LeftShift(Quire,Int32).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := AfterFinished;
                                    \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= true;
                                    \Quire Quire::op_LeftShift(Quire,Int32).0._Started\ <= false;
                                    \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).return.0\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.return\;
                                    \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32).left.parameter.In.0\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.left.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire Quire::op_LeftShift(Quire,Int32).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForStarted;
                            \Quire Posit32::op_Explicit(Posit32).0.Quire Quire::op_LeftShift(Quire,Int32)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    


    
    
    \UInt32 Quire::op_Explicit(Quire).0._Started\ <= \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire)._Started.0\;
    \UInt32 Quire::op_Explicit(Quire).0.x.parameter.In\ <= \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire).x.parameter.Out.0\;
    \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire)._Finished.0\ <= \UInt32 Quire::op_Explicit(Quire).0._Finished\;
    \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire).return.0\ <= \UInt32 Quire::op_Explicit(Quire).0.return\;
    \Posit32::.ctor(Quire).0.UInt32 Quire::op_Explicit(Quire).x.parameter.In.0\ <= \UInt32 Quire::op_Explicit(Quire).0.x.parameter.Out\;
    


    
    
    \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._Started\ <= \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32)._Started.0\;
    \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.signBit.parameter.In\ <= \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).signBit.parameter.Out.0\;
    \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.regimeKValue.parameter.In\ <= \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).regimeKValue.parameter.Out.0\;
    \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.exponentBits.parameter.In\ <= \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).exponentBits.parameter.Out.0\;
    \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.fractionBits.parameter.In\ <= \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).fractionBits.parameter.Out.0\;
    \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32)._Finished.0\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0._Finished\;
    \Posit32::.ctor(Quire).0.Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).return.0\ <= \Posit32::AssemblePositBitsWithRounding(Boolean,Int32,UInt32,UInt32).0.return\;
    


    
    
    \Posit32::.ctor(UInt32).0._Started\ <= \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32)._Started.0\;
    \Posit32::.ctor(UInt32).0.this.parameter.In\ <= \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32).this.parameter.Out.0\;
    \Posit32::.ctor(UInt32).0.value.parameter.In\ <= \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32).value.parameter.Out.0\;
    \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32)._Finished.0\ <= \Posit32::.ctor(UInt32).0._Finished\;
    \Posit32::.ctor(Int32).0.Posit32::.ctor(UInt32).this.parameter.In.0\ <= \Posit32::.ctor(UInt32).0.this.parameter.Out\;
    


    
    \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Posit32::op_Explicit(Posit32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Quire::op_Addition(Quire,UInt32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Quire::op_Addition(Quire,UInt32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\ := WaitingForStarted;
                \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Finished.0\ <= false;
                \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16)._Finished.0\ <= false;
                \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Finished.0\ <= false;
            else 

                
                case \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Started.0\) then 
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ := 0;
                            \Quire::.ctor(UInt32,UInt16).0._Started\ <= true;
                            \Quire::.ctor(UInt32,UInt16).0.this.parameter.In\ <= \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).this.parameter.Out.0\;
                            \Quire::.ctor(UInt32,UInt16).0.firstSegment.parameter.In\ <= \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).firstSegment.parameter.Out.0\;
                            \Quire::.ctor(UInt32,UInt16).0.size.parameter.In\ <= \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire::.ctor(UInt32,UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := AfterFinished;
                                    \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Finished.0\ <= true;
                                    \Quire::.ctor(UInt32,UInt16).0._Started\ <= false;
                                    \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16).this.parameter.In.0\ <= \Quire::.ctor(UInt32,UInt16).0.this.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForStarted;
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire::.ctor(UInt32,UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16)._Started.0\) then 
                            \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ := 0;
                            \Quire::.ctor(UInt32,UInt16).0._Started\ <= true;
                            \Quire::.ctor(UInt32,UInt16).0.this.parameter.In\ <= \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16).this.parameter.Out.0\;
                            \Quire::.ctor(UInt32,UInt16).0.firstSegment.parameter.In\ <= \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16).firstSegment.parameter.Out.0\;
                            \Quire::.ctor(UInt32,UInt16).0.size.parameter.In\ <= \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire::.ctor(UInt32,UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := AfterFinished;
                                    \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16)._Finished.0\ <= true;
                                    \Quire::.ctor(UInt32,UInt16).0._Started\ <= false;
                                    \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16).this.parameter.In.0\ <= \Quire::.ctor(UInt32,UInt16).0.this.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForStarted;
                            \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt32,UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Started.0\) then 
                            \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Quire::op_Addition(Quire,UInt32).0.runningIndex.0\ := 0;
                            \Quire::.ctor(UInt32,UInt16).0._Started\ <= true;
                            \Quire::.ctor(UInt32,UInt16).0.this.parameter.In\ <= \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).this.parameter.Out.0\;
                            \Quire::.ctor(UInt32,UInt16).0.firstSegment.parameter.In\ <= \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).firstSegment.parameter.Out.0\;
                            \Quire::.ctor(UInt32,UInt16).0.size.parameter.In\ <= \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Quire::op_Addition(Quire,UInt32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire::.ctor(UInt32,UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\ := AfterFinished;
                                    \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Finished.0\ <= true;
                                    \Quire::.ctor(UInt32,UInt16).0._Started\ <= false;
                                    \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16).this.parameter.In.0\ <= \Quire::.ctor(UInt32,UInt16).0.this.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt32,UInt16).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\ := WaitingForStarted;
                            \Quire Quire::op_Addition(Quire,UInt32).0.Quire::.ctor(UInt32,UInt16)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    


    
    
    \Boolean Quire::op_Equality(Quire,Quire).0._Started\ <= \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire)._Started.0\;
    \Boolean Quire::op_Equality(Quire,Quire).0.left.parameter.In\ <= \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).left.parameter.Out.0\;
    \Boolean Quire::op_Equality(Quire,Quire).0.right.parameter.In\ <= \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).right.parameter.Out.0\;
    \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire)._Finished.0\ <= \Boolean Quire::op_Equality(Quire,Quire).0._Finished\;
    \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).return.0\ <= \Boolean Quire::op_Equality(Quire,Quire).0.return\;
    \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).left.parameter.In.0\ <= \Boolean Quire::op_Equality(Quire,Quire).0.left.parameter.Out\;
    \Posit32::FusedSum(Posit32[],Quire).0.Boolean Quire::op_Equality(Quire,Quire).right.parameter.In.0\ <= \Boolean Quire::op_Equality(Quire,Quire).0.right.parameter.Out\;
    


    
    \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Quire Quire::op_Addition(Quire,UInt32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Quire Quire::op_Addition(Quire,UInt32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\ := WaitingForStarted;
                \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\ <= false;
                \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\ <= false;
            else 

                
                case \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\) then 
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ := 0;
                            \Quire Quire::op_Addition(Quire,Quire).0._Started\ <= true;
                            \Quire Quire::op_Addition(Quire,Quire).0.left.parameter.In\ <= \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.Out.0\;
                            \Quire Quire::op_Addition(Quire,Quire).0.right.parameter.In\ <= \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Posit32::FusedSum(Posit32[],Quire).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire Quire::op_Addition(Quire,Quire).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := AfterFinished;
                                    \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\ <= true;
                                    \Quire Quire::op_Addition(Quire,Quire).0._Started\ <= false;
                                    \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).return.0\ <= \Quire Quire::op_Addition(Quire,Quire).0.return\;
                                    \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.In.0\ <= \Quire Quire::op_Addition(Quire,Quire).0.left.parameter.Out\;
                                    \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.In.0\ <= \Quire Quire::op_Addition(Quire,Quire).0.right.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Posit32::FusedSum(Posit32[],Quire).0.runningState.0\ := WaitingForStarted;
                            \Posit32::FusedSum(Posit32[],Quire).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\) then 
                            \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Quire Quire::op_Addition(Quire,UInt32).0.runningIndex.0\ := 0;
                            \Quire Quire::op_Addition(Quire,Quire).0._Started\ <= true;
                            \Quire Quire::op_Addition(Quire,Quire).0.left.parameter.In\ <= \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.Out.0\;
                            \Quire Quire::op_Addition(Quire,Quire).0.right.parameter.In\ <= \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Quire Quire::op_Addition(Quire,UInt32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire Quire::op_Addition(Quire,Quire).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\ := AfterFinished;
                                    \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\ <= true;
                                    \Quire Quire::op_Addition(Quire,Quire).0._Started\ <= false;
                                    \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).return.0\ <= \Quire Quire::op_Addition(Quire,Quire).0.return\;
                                    \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).left.parameter.In.0\ <= \Quire Quire::op_Addition(Quire,Quire).0.left.parameter.Out\;
                                    \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire).right.parameter.In.0\ <= \Quire Quire::op_Addition(Quire,Quire).0.right.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire Quire::op_Addition(Quire,Quire).Quire Quire::op_Addition(Quire,UInt32).0.runningState.0\ := WaitingForStarted;
                            \Quire Quire::op_Addition(Quire,UInt32).0.Quire Quire::op_Addition(Quire,Quire)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    


    
    \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16)\: process (\Clock\) 
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Posit32::op_Explicit(Posit32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_Addition(Quire,Quire).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_Addition(Quire,Quire).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_RightShift(Quire,Int32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_RightShift(Quire,Int32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_LeftShift(Quire,Int32).0.runningIndex.0\: integer range 0 to 0 := 0;
        Variable \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_LeftShift(Quire,Int32).0.runningState.0\: \Hast::InternalInvocationProxy()._RunningStates\ := WaitingForStarted;
    begin 
        if (rising_edge(\Clock\)) then 
            if (\Reset\ = '1') then 
                
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_Addition(Quire,Quire).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_Addition(Quire,Quire).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_RightShift(Quire,Int32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_RightShift(Quire,Int32).0.runningState.0\ := WaitingForStarted;
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_LeftShift(Quire,Int32).0.runningIndex.0\ := 0;
                \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_LeftShift(Quire,Int32).0.runningState.0\ := WaitingForStarted;
                \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
                \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
                \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
                \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
            else 

                
                case \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\) then 
                            \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ := 0;
                            \Quire::.ctor(UInt64[],UInt16).0._Started\ <= true;
                            \Quire::.ctor(UInt64[],UInt16).0.this.parameter.In\ <= \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\;
                            \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.In\ <= \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\;
                            \Quire::.ctor(UInt64[],UInt16).0.size.parameter.In\ <= \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Posit32::op_Explicit(Posit32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire::.ctor(UInt64[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := AfterFinished;
                                    \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= true;
                                    \Quire::.ctor(UInt64[],UInt16).0._Started\ <= false;
                                    \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\ <= \Quire::.ctor(UInt64[],UInt16).0.this.parameter.Out\;
                                    \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\ <= \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Posit32::op_Explicit(Posit32).0.runningState.0\ := WaitingForStarted;
                            \Quire Posit32::op_Explicit(Posit32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_Addition(Quire,Quire).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Started.0\) then 
                            \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_Addition(Quire,Quire).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_Addition(Quire,Quire).0.runningIndex.0\ := 0;
                            \Quire::.ctor(UInt64[],UInt16).0._Started\ <= true;
                            \Quire::.ctor(UInt64[],UInt16).0.this.parameter.In\ <= \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\;
                            \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.In\ <= \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\;
                            \Quire::.ctor(UInt64[],UInt16).0.size.parameter.In\ <= \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_Addition(Quire,Quire).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire::.ctor(UInt64[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_Addition(Quire,Quire).0.runningState.0\ := AfterFinished;
                                    \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= true;
                                    \Quire::.ctor(UInt64[],UInt16).0._Started\ <= false;
                                    \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\ <= \Quire::.ctor(UInt64[],UInt16).0.this.parameter.Out\;
                                    \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\ <= \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_Addition(Quire,Quire).0.runningState.0\ := WaitingForStarted;
                            \Quire Quire::op_Addition(Quire,Quire).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_RightShift(Quire,Int32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\) then 
                            \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_RightShift(Quire,Int32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_RightShift(Quire,Int32).0.runningIndex.0\ := 0;
                            \Quire::.ctor(UInt64[],UInt16).0._Started\ <= true;
                            \Quire::.ctor(UInt64[],UInt16).0.this.parameter.In\ <= \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\;
                            \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.In\ <= \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\;
                            \Quire::.ctor(UInt64[],UInt16).0.size.parameter.In\ <= \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_RightShift(Quire,Int32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire::.ctor(UInt64[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_RightShift(Quire,Int32).0.runningState.0\ := AfterFinished;
                                    \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= true;
                                    \Quire::.ctor(UInt64[],UInt16).0._Started\ <= false;
                                    \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\ <= \Quire::.ctor(UInt64[],UInt16).0.this.parameter.Out\;
                                    \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\ <= \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_RightShift(Quire,Int32).0.runningState.0\ := WaitingForStarted;
                            \Quire Quire::op_RightShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;


                
                case \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_LeftShift(Quire,Int32).0.runningState.0\ is 
                    when WaitingForStarted => 
                        if (\Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\) then 
                            \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_LeftShift(Quire,Int32).0.runningState.0\ := WaitingForFinished;
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_LeftShift(Quire,Int32).0.runningIndex.0\ := 0;
                            \Quire::.ctor(UInt64[],UInt16).0._Started\ <= true;
                            \Quire::.ctor(UInt64[],UInt16).0.this.parameter.In\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.Out.0\;
                            \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.In\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.Out.0\;
                            \Quire::.ctor(UInt64[],UInt16).0.size.parameter.In\ <= \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).size.parameter.Out.0\;
                        end if;
                    when WaitingForFinished => 
                        case \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_LeftShift(Quire,Int32).0.runningIndex.0\ is 
                            when 0 => 
                                if (\Quire::.ctor(UInt64[],UInt16).0._Finished\) then 
                                    \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_LeftShift(Quire,Int32).0.runningState.0\ := AfterFinished;
                                    \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= true;
                                    \Quire::.ctor(UInt64[],UInt16).0._Started\ <= false;
                                    \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).this.parameter.In.0\ <= \Quire::.ctor(UInt64[],UInt16).0.this.parameter.Out\;
                                    \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16).segments.parameter.In.0\ <= \Quire::.ctor(UInt64[],UInt16).0.segments.parameter.Out\;
                                end if;
                        end case;
                    when AfterFinished => 
                        
                        if (\Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Started.0\ = false) then 
                            \Hast::InternalInvocationProxy().Quire::.ctor(UInt64[],UInt16).Quire Quire::op_LeftShift(Quire,Int32).0.runningState.0\ := WaitingForStarted;
                            \Quire Quire::op_LeftShift(Quire,Int32).0.Quire::.ctor(UInt64[],UInt16)._Finished.0\ <= false;
                        end if;
                end case;

            end if;
        end if;
    end process;
    


    
    
    \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._Started\ <= \Hast::ExternalInvocationProxy().Posit32FusedCalculator::CalculateFusedSum(SimpleMemory)._Started.0\;
    \Hast::ExternalInvocationProxy().Posit32FusedCalculator::CalculateFusedSum(SimpleMemory)._Finished.0\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0._Finished\;
    


    
    \CellIndex\ <= to_integer(\Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.CellIndex\) when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.ReadEnable\ or \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.WriteEnable\ else 0;
    \DataOut\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.DataOut\ when \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.WriteEnable\ else (others => '0');
    \ReadEnable\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.ReadEnable\;
    \WriteEnable\ <= \Posit32FusedCalculator::CalculateFusedSum(SimpleMemory).0.SimpleMemory.WriteEnable\;
    

end Imp;
